`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/16/2023 08:13:15 PM
// Design Name: 
// Module Name: leg_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module leg_rom(
    input clk_i,
    input [11:0] addr,
    output reg [11:0] color_o
    );

reg[11:0] addr_in;

always @ (posedge clk_i) begin
    addr_in <= addr;            // latch in current address
end    
    
always @*
    case(addr_in)
		12'd0: color_o = 12'b000011110000;
		12'd1: color_o = 12'b000000000000;
		12'd2: color_o = 12'b000000000000;
		12'd3: color_o = 12'b000000000000;
		12'd4: color_o = 12'b000000000000;
		12'd5: color_o = 12'b100000000001;
		12'd6: color_o = 12'b100000000001;
		12'd7: color_o = 12'b100000000001;
		12'd8: color_o = 12'b100000000001;
		12'd9: color_o = 12'b000000000000;
		12'd10: color_o = 12'b000000000000;
		12'd11: color_o = 12'b000000000000;
		12'd12: color_o = 12'b000000000000;
		12'd13: color_o = 12'b000000000000;
		12'd14: color_o = 12'b100000000000;
		12'd15: color_o = 12'b100000000000;
		12'd16: color_o = 12'b100000000000;
		12'd17: color_o = 12'b100000000000;
		12'd18: color_o = 12'b000000000000;
		12'd19: color_o = 12'b100000000000;
		12'd20: color_o = 12'b100000000001;
		12'd21: color_o = 12'b100000000001;
		12'd22: color_o = 12'b000000000000;
		12'd23: color_o = 12'b000011110000;
		12'd24: color_o = 12'b000011110000;
		12'd25: color_o = 12'b000011110000;
		12'd26: color_o = 12'b000011110000;
		12'd27: color_o = 12'b000011110000;
		12'd28: color_o = 12'b000011110000;
		12'd29: color_o = 12'b000011110000;
		12'd30: color_o = 12'b000011110000;
		12'd31: color_o = 12'b000011110000;
		12'd32: color_o = 12'b000011110000;
		12'd33: color_o = 12'b000000000000;
		12'd34: color_o = 12'b000000000000;
		12'd35: color_o = 12'b000000000000;
		12'd36: color_o = 12'b000000000000;
		12'd37: color_o = 12'b000000000000;
		12'd38: color_o = 12'b000000000000;
		12'd39: color_o = 12'b100000000000;
		12'd40: color_o = 12'b100000000001;
		12'd41: color_o = 12'b100000000001;
		12'd42: color_o = 12'b100000000000;
		12'd43: color_o = 12'b100000000000;
		12'd44: color_o = 12'b100000000000;
		12'd45: color_o = 12'b100000000000;
		12'd46: color_o = 12'b010000000000;
		12'd47: color_o = 12'b010000000000;
		12'd48: color_o = 12'b010000000000;
		12'd49: color_o = 12'b010000000000;
		12'd50: color_o = 12'b000000000000;
		12'd51: color_o = 12'b000000000000;
		12'd52: color_o = 12'b000000000000;
		12'd53: color_o = 12'b100000000001;
		12'd54: color_o = 12'b000000000000;
		12'd55: color_o = 12'b000011110000;
		12'd56: color_o = 12'b000011110000;
		12'd57: color_o = 12'b000011110000;
		12'd58: color_o = 12'b000011110000;
		12'd59: color_o = 12'b000011110000;
		12'd60: color_o = 12'b000011110000;
		12'd61: color_o = 12'b000011110000;
		12'd62: color_o = 12'b000011110000;
		12'd63: color_o = 12'b000011110000;
		12'd64: color_o = 12'b000011110000;
		12'd65: color_o = 12'b000000000000;
		12'd66: color_o = 12'b000000000000;
		12'd67: color_o = 12'b000000000000;
		12'd68: color_o = 12'b100000000001;
		12'd69: color_o = 12'b100000000001;
		12'd70: color_o = 12'b000000000000;
		12'd71: color_o = 12'b000000000000;
		12'd72: color_o = 12'b000000000000;
		12'd73: color_o = 12'b000000000000;
		12'd74: color_o = 12'b100000000000;
		12'd75: color_o = 12'b010000000000;
		12'd76: color_o = 12'b010000000000;
		12'd77: color_o = 12'b010000000000;
		12'd78: color_o = 12'b010000000000;
		12'd79: color_o = 12'b010000000000;
		12'd80: color_o = 12'b000000000000;
		12'd81: color_o = 12'b000000000000;
		12'd82: color_o = 12'b000000000000;
		12'd83: color_o = 12'b010000000000;
		12'd84: color_o = 12'b010000000000;
		12'd85: color_o = 12'b000000000000;
		12'd86: color_o = 12'b000000000000;
		12'd87: color_o = 12'b000011110000;
		12'd88: color_o = 12'b000011110000;
		12'd89: color_o = 12'b000011110000;
		12'd90: color_o = 12'b000011110000;
		12'd91: color_o = 12'b000011110000;
		12'd92: color_o = 12'b000011110000;
		12'd93: color_o = 12'b000011110000;
		12'd94: color_o = 12'b000011110000;
		12'd95: color_o = 12'b000011110000;
		12'd96: color_o = 12'b000011110000;
		12'd97: color_o = 12'b000011110000;
		12'd98: color_o = 12'b000000000000;
		12'd99: color_o = 12'b000000000000;
		12'd100: color_o = 12'b100000000001;
		12'd101: color_o = 12'b000000000000;
		12'd102: color_o = 12'b000000000000;
		12'd103: color_o = 12'b000000000000;
		12'd104: color_o = 12'b000000000000;
		12'd105: color_o = 12'b000000000000;
		12'd106: color_o = 12'b000000000000;
		12'd107: color_o = 12'b000000000000;
		12'd108: color_o = 12'b000000000000;
		12'd109: color_o = 12'b000000000000;
		12'd110: color_o = 12'b000000000000;
		12'd111: color_o = 12'b000000000000;
		12'd112: color_o = 12'b000000000000;
		12'd113: color_o = 12'b000000000000;
		12'd114: color_o = 12'b100000000001;
		12'd115: color_o = 12'b100000000001;
		12'd116: color_o = 12'b000000000000;
		12'd117: color_o = 12'b000000000000;
		12'd118: color_o = 12'b000011110000;
		12'd119: color_o = 12'b000011110000;
		12'd120: color_o = 12'b000011110000;
		12'd121: color_o = 12'b000011110000;
		12'd122: color_o = 12'b000011110000;
		12'd123: color_o = 12'b000011110000;
		12'd124: color_o = 12'b000011110000;
		12'd125: color_o = 12'b000011110000;
		12'd126: color_o = 12'b000011110000;
		12'd127: color_o = 12'b000011110000;
		12'd128: color_o = 12'b000011110000;
		12'd129: color_o = 12'b000011110000;
		12'd130: color_o = 12'b000000000000;
		12'd131: color_o = 12'b100000000001;
		12'd132: color_o = 12'b100000000001;
		12'd133: color_o = 12'b100000000001;
		12'd134: color_o = 12'b100000000001;
		12'd135: color_o = 12'b100000000001;
		12'd136: color_o = 12'b010000000000;
		12'd137: color_o = 12'b100000000001;
		12'd138: color_o = 12'b100000000001;
		12'd139: color_o = 12'b100000000001;
		12'd140: color_o = 12'b100000000001;
		12'd141: color_o = 12'b100000000001;
		12'd142: color_o = 12'b100000000001;
		12'd143: color_o = 12'b100000000001;
		12'd144: color_o = 12'b100000000001;
		12'd145: color_o = 12'b100000000001;
		12'd146: color_o = 12'b100000000001;
		12'd147: color_o = 12'b100000000001;
		12'd148: color_o = 12'b000000000000;
		12'd149: color_o = 12'b000011110000;
		12'd150: color_o = 12'b000011110000;
		12'd151: color_o = 12'b000011110000;
		12'd152: color_o = 12'b000011110000;
		12'd153: color_o = 12'b000011110000;
		12'd154: color_o = 12'b000011110000;
		12'd155: color_o = 12'b000011110000;
		12'd156: color_o = 12'b000011110000;
		12'd157: color_o = 12'b000011110000;
		12'd158: color_o = 12'b000011110000;
		12'd159: color_o = 12'b000011110000;
		12'd160: color_o = 12'b000011110000;
		12'd161: color_o = 12'b000011110000;
		12'd162: color_o = 12'b000000000000;
		12'd163: color_o = 12'b000000000000;
		12'd164: color_o = 12'b100000000001;
		12'd165: color_o = 12'b100000000001;
		12'd166: color_o = 12'b010000000000;
		12'd167: color_o = 12'b010000000000;
		12'd168: color_o = 12'b100000000001;
		12'd169: color_o = 12'b010000000000;
		12'd170: color_o = 12'b100000000001;
		12'd171: color_o = 12'b100000000001;
		12'd172: color_o = 12'b100000000001;
		12'd173: color_o = 12'b100000000001;
		12'd174: color_o = 12'b100000000001;
		12'd175: color_o = 12'b100000000001;
		12'd176: color_o = 12'b100000000001;
		12'd177: color_o = 12'b100000000001;
		12'd178: color_o = 12'b100000000001;
		12'd179: color_o = 12'b100000000001;
		12'd180: color_o = 12'b000000000000;
		12'd181: color_o = 12'b000011110000;
		12'd182: color_o = 12'b000011110000;
		12'd183: color_o = 12'b000011110000;
		12'd184: color_o = 12'b000011110000;
		12'd185: color_o = 12'b000011110000;
		12'd186: color_o = 12'b000011110000;
		12'd187: color_o = 12'b000011110000;
		12'd188: color_o = 12'b000011110000;
		12'd189: color_o = 12'b000011110000;
		12'd190: color_o = 12'b000011110000;
		12'd191: color_o = 12'b000011110000;
		12'd192: color_o = 12'b000011110000;
		12'd193: color_o = 12'b000011110000;
		12'd194: color_o = 12'b000000000000;
		12'd195: color_o = 12'b000000000000;
		12'd196: color_o = 12'b100000000001;
		12'd197: color_o = 12'b000000000000;
		12'd198: color_o = 12'b010000000000;
		12'd199: color_o = 12'b100000000001;
		12'd200: color_o = 12'b010000000000;
		12'd201: color_o = 12'b100000000001;
		12'd202: color_o = 12'b100000000001;
		12'd203: color_o = 12'b100000000001;
		12'd204: color_o = 12'b100000000001;
		12'd205: color_o = 12'b100000000001;
		12'd206: color_o = 12'b100000000001;
		12'd207: color_o = 12'b000000000000;
		12'd208: color_o = 12'b000000000000;
		12'd209: color_o = 12'b100000000001;
		12'd210: color_o = 12'b100000000001;
		12'd211: color_o = 12'b000000000000;
		12'd212: color_o = 12'b000011110000;
		12'd213: color_o = 12'b000011110000;
		12'd214: color_o = 12'b000011110000;
		12'd215: color_o = 12'b000011110000;
		12'd216: color_o = 12'b000011110000;
		12'd217: color_o = 12'b000011110000;
		12'd218: color_o = 12'b000011110000;
		12'd219: color_o = 12'b000011110000;
		12'd220: color_o = 12'b000011110000;
		12'd221: color_o = 12'b000011110000;
		12'd222: color_o = 12'b000011110000;
		12'd223: color_o = 12'b000011110000;
		12'd224: color_o = 12'b000011110000;
		12'd225: color_o = 12'b000011110000;
		12'd226: color_o = 12'b000011110000;
		12'd227: color_o = 12'b000000000000;
		12'd228: color_o = 12'b000000000000;
		12'd229: color_o = 12'b000000000000;
		12'd230: color_o = 12'b010000000000;
		12'd231: color_o = 12'b010000000000;
		12'd232: color_o = 12'b100000000001;
		12'd233: color_o = 12'b100000000001;
		12'd234: color_o = 12'b100000000001;
		12'd235: color_o = 12'b100000000001;
		12'd236: color_o = 12'b100000000001;
		12'd237: color_o = 12'b100000000001;
		12'd238: color_o = 12'b000000000000;
		12'd239: color_o = 12'b000000000000;
		12'd240: color_o = 12'b010000000000;
		12'd241: color_o = 12'b100000000001;
		12'd242: color_o = 12'b000000000000;
		12'd243: color_o = 12'b000011110000;
		12'd244: color_o = 12'b000011110000;
		12'd245: color_o = 12'b000011110000;
		12'd246: color_o = 12'b000011110000;
		12'd247: color_o = 12'b000011110000;
		12'd248: color_o = 12'b000011110000;
		12'd249: color_o = 12'b000011110000;
		12'd250: color_o = 12'b000011110000;
		12'd251: color_o = 12'b000011110000;
		12'd252: color_o = 12'b000011110000;
		12'd253: color_o = 12'b000011110000;
		12'd254: color_o = 12'b000011110000;
		12'd255: color_o = 12'b000011110000;
		12'd256: color_o = 12'b000011110000;
		12'd257: color_o = 12'b000011110000;
		12'd258: color_o = 12'b000011110000;
		12'd259: color_o = 12'b000011110000;
		12'd260: color_o = 12'b000000000000;
		12'd261: color_o = 12'b000000000000;
		12'd262: color_o = 12'b010000000000;
		12'd263: color_o = 12'b100000000001;
		12'd264: color_o = 12'b100000000001;
		12'd265: color_o = 12'b100000000001;
		12'd266: color_o = 12'b100000000001;
		12'd267: color_o = 12'b100000000001;
		12'd268: color_o = 12'b100000000001;
		12'd269: color_o = 12'b100000000001;
		12'd270: color_o = 12'b000000000000;
		12'd271: color_o = 12'b010000000000;
		12'd272: color_o = 12'b100000000001;
		12'd273: color_o = 12'b000000000000;
		12'd274: color_o = 12'b000000000000;
		12'd275: color_o = 12'b000011110000;
		12'd276: color_o = 12'b000011110000;
		12'd277: color_o = 12'b000011110000;
		12'd278: color_o = 12'b000011110000;
		12'd279: color_o = 12'b000011110000;
		12'd280: color_o = 12'b000011110000;
		12'd281: color_o = 12'b000011110000;
		12'd282: color_o = 12'b000011110000;
		12'd283: color_o = 12'b000011110000;
		12'd284: color_o = 12'b000011110000;
		12'd285: color_o = 12'b000011110000;
		12'd286: color_o = 12'b000011110000;
		12'd287: color_o = 12'b000011110000;
		12'd288: color_o = 12'b000011110000;
		12'd289: color_o = 12'b000011110000;
		12'd290: color_o = 12'b000011110000;
		12'd291: color_o = 12'b000011110000;
		12'd292: color_o = 12'b000011110000;
		12'd293: color_o = 12'b000000000000;
		12'd294: color_o = 12'b010000000000;
		12'd295: color_o = 12'b010000000000;
		12'd296: color_o = 12'b100000000001;
		12'd297: color_o = 12'b010000000000;
		12'd298: color_o = 12'b100000000001;
		12'd299: color_o = 12'b100000000001;
		12'd300: color_o = 12'b100000000001;
		12'd301: color_o = 12'b000000000000;
		12'd302: color_o = 12'b000000000000;
		12'd303: color_o = 12'b100000000001;
		12'd304: color_o = 12'b010000000000;
		12'd305: color_o = 12'b100000000001;
		12'd306: color_o = 12'b000000000000;
		12'd307: color_o = 12'b000011110000;
		12'd308: color_o = 12'b000011110000;
		12'd309: color_o = 12'b000011110000;
		12'd310: color_o = 12'b000011110000;
		12'd311: color_o = 12'b000011110000;
		12'd312: color_o = 12'b000011110000;
		12'd313: color_o = 12'b000011110000;
		12'd314: color_o = 12'b000011110000;
		12'd315: color_o = 12'b000011110000;
		12'd316: color_o = 12'b000011110000;
		12'd317: color_o = 12'b000011110000;
		12'd318: color_o = 12'b000011110000;
		12'd319: color_o = 12'b000011110000;
		12'd320: color_o = 12'b000011110000;
		12'd321: color_o = 12'b000011110000;
		12'd322: color_o = 12'b000011110000;
		12'd323: color_o = 12'b000011110000;
		12'd324: color_o = 12'b000011110000;
		12'd325: color_o = 12'b000011110000;
		12'd326: color_o = 12'b000000000000;
		12'd327: color_o = 12'b010000000000;
		12'd328: color_o = 12'b010000000000;
		12'd329: color_o = 12'b010000000000;
		12'd330: color_o = 12'b100000000001;
		12'd331: color_o = 12'b100000000001;
		12'd332: color_o = 12'b100000000001;
		12'd333: color_o = 12'b000000000000;
		12'd334: color_o = 12'b100000000001;
		12'd335: color_o = 12'b010000000000;
		12'd336: color_o = 12'b100000000001;
		12'd337: color_o = 12'b000000000000;
		12'd338: color_o = 12'b000011110000;
		12'd339: color_o = 12'b000011110000;
		12'd340: color_o = 12'b000011110000;
		12'd341: color_o = 12'b000011110000;
		12'd342: color_o = 12'b000011110000;
		12'd343: color_o = 12'b000011110000;
		12'd344: color_o = 12'b000011110000;
		12'd345: color_o = 12'b000011110000;
		12'd346: color_o = 12'b000011110000;
		12'd347: color_o = 12'b000011110000;
		12'd348: color_o = 12'b000011110000;
		12'd349: color_o = 12'b000011110000;
		12'd350: color_o = 12'b000011110000;
		12'd351: color_o = 12'b000011110000;
		12'd352: color_o = 12'b000011110000;
		12'd353: color_o = 12'b000011110000;
		12'd354: color_o = 12'b000011110000;
		12'd355: color_o = 12'b000011110000;
		12'd356: color_o = 12'b000011110000;
		12'd357: color_o = 12'b000011110000;
		12'd358: color_o = 12'b000000000000;
		12'd359: color_o = 12'b010000000000;
		12'd360: color_o = 12'b010000000000;
		12'd361: color_o = 12'b100000000001;
		12'd362: color_o = 12'b010000000000;
		12'd363: color_o = 12'b100000000001;
		12'd364: color_o = 12'b100000000001;
		12'd365: color_o = 12'b100000000001;
		12'd366: color_o = 12'b100000000001;
		12'd367: color_o = 12'b000000000000;
		12'd368: color_o = 12'b000000000000;
		12'd369: color_o = 12'b000000000000;
		12'd370: color_o = 12'b000011110000;
		12'd371: color_o = 12'b000011110000;
		12'd372: color_o = 12'b000011110000;
		12'd373: color_o = 12'b000011110000;
		12'd374: color_o = 12'b000011110000;
		12'd375: color_o = 12'b000011110000;
		12'd376: color_o = 12'b000011110000;
		12'd377: color_o = 12'b000011110000;
		12'd378: color_o = 12'b000011110000;
		12'd379: color_o = 12'b000011110000;
		12'd380: color_o = 12'b000011110000;
		12'd381: color_o = 12'b000011110000;
		12'd382: color_o = 12'b000011110000;
		12'd383: color_o = 12'b000011110000;
		12'd384: color_o = 12'b000011110000;
		12'd385: color_o = 12'b000011110000;
		12'd386: color_o = 12'b000011110000;
		12'd387: color_o = 12'b000011110000;
		12'd388: color_o = 12'b000011110000;
		12'd389: color_o = 12'b000011110000;
		12'd390: color_o = 12'b000000000000;
		12'd391: color_o = 12'b010000000000;
		12'd392: color_o = 12'b010000000000;
		12'd393: color_o = 12'b010000000000;
		12'd394: color_o = 12'b100000000001;
		12'd395: color_o = 12'b100000000001;
		12'd396: color_o = 12'b100000000001;
		12'd397: color_o = 12'b100000000001;
		12'd398: color_o = 12'b100000000001;
		12'd399: color_o = 12'b010000000000;
		12'd400: color_o = 12'b000000000000;
		12'd401: color_o = 12'b000011110000;
		12'd402: color_o = 12'b000011110000;
		12'd403: color_o = 12'b000011110000;
		12'd404: color_o = 12'b000011110000;
		12'd405: color_o = 12'b000011110000;
		12'd406: color_o = 12'b000011110000;
		12'd407: color_o = 12'b000011110000;
		12'd408: color_o = 12'b000011110000;
		12'd409: color_o = 12'b000011110000;
		12'd410: color_o = 12'b000011110000;
		12'd411: color_o = 12'b000011110000;
		12'd412: color_o = 12'b000011110000;
		12'd413: color_o = 12'b000011110000;
		12'd414: color_o = 12'b000011110000;
		12'd415: color_o = 12'b000011110000;
		12'd416: color_o = 12'b000011110000;
		12'd417: color_o = 12'b000011110000;
		12'd418: color_o = 12'b000011110000;
		12'd419: color_o = 12'b000011110000;
		12'd420: color_o = 12'b000011110000;
		12'd421: color_o = 12'b000011110000;
		12'd422: color_o = 12'b000000000000;
		12'd423: color_o = 12'b000000000000;
		12'd424: color_o = 12'b000000000000;
		12'd425: color_o = 12'b100000000001;
		12'd426: color_o = 12'b010000000000;
		12'd427: color_o = 12'b100000000001;
		12'd428: color_o = 12'b100000000001;
		12'd429: color_o = 12'b100000000001;
		12'd430: color_o = 12'b100000000001;
		12'd431: color_o = 12'b100000000001;
		12'd432: color_o = 12'b000000000000;
		12'd433: color_o = 12'b000000000000;
		12'd434: color_o = 12'b000011110000;
		12'd435: color_o = 12'b000011110000;
		12'd436: color_o = 12'b000011110000;
		12'd437: color_o = 12'b000011110000;
		12'd438: color_o = 12'b000011110000;
		12'd439: color_o = 12'b000011110000;
		12'd440: color_o = 12'b000011110000;
		12'd441: color_o = 12'b000011110000;
		12'd442: color_o = 12'b000011110000;
		12'd443: color_o = 12'b000011110000;
		12'd444: color_o = 12'b000011110000;
		12'd445: color_o = 12'b000011110000;
		12'd446: color_o = 12'b000011110000;
		12'd447: color_o = 12'b000011110000;
		12'd448: color_o = 12'b000011110000;
		12'd449: color_o = 12'b000011110000;
		12'd450: color_o = 12'b000011110000;
		12'd451: color_o = 12'b000011110000;
		12'd452: color_o = 12'b000011110000;
		12'd453: color_o = 12'b000011110000;
		12'd454: color_o = 12'b000011110000;
		12'd455: color_o = 12'b000000000000;
		12'd456: color_o = 12'b000000000000;
		12'd457: color_o = 12'b010000000000;
		12'd458: color_o = 12'b100000000001;
		12'd459: color_o = 12'b010000000000;
		12'd460: color_o = 12'b100000000001;
		12'd461: color_o = 12'b100000000001;
		12'd462: color_o = 12'b100000000001;
		12'd463: color_o = 12'b000000000000;
		12'd464: color_o = 12'b000000000000;
		12'd465: color_o = 12'b000000000000;
		12'd466: color_o = 12'b000000000000;
		12'd467: color_o = 12'b000011110000;
		12'd468: color_o = 12'b000011110000;
		12'd469: color_o = 12'b000011110000;
		12'd470: color_o = 12'b000011110000;
		12'd471: color_o = 12'b000011110000;
		12'd472: color_o = 12'b000011110000;
		12'd473: color_o = 12'b000011110000;
		12'd474: color_o = 12'b000011110000;
		12'd475: color_o = 12'b000011110000;
		12'd476: color_o = 12'b000011110000;
		12'd477: color_o = 12'b000011110000;
		12'd478: color_o = 12'b000011110000;
		12'd479: color_o = 12'b000011110000;
		12'd480: color_o = 12'b000011110000;
		12'd481: color_o = 12'b000011110000;
		12'd482: color_o = 12'b000011110000;
		12'd483: color_o = 12'b000011110000;
		12'd484: color_o = 12'b000011110000;
		12'd485: color_o = 12'b000011110000;
		12'd486: color_o = 12'b000011110000;
		12'd487: color_o = 12'b000011110000;
		12'd488: color_o = 12'b000000000000;
		12'd489: color_o = 12'b000000000000;
		12'd490: color_o = 12'b000000000000;
		12'd491: color_o = 12'b100000000001;
		12'd492: color_o = 12'b010000000000;
		12'd493: color_o = 12'b100000000001;
		12'd494: color_o = 12'b000000000000;
		12'd495: color_o = 12'b000000000000;
		12'd496: color_o = 12'b000000000000;
		12'd497: color_o = 12'b000000000000;
		12'd498: color_o = 12'b000000000000;
		12'd499: color_o = 12'b000000000000;
		12'd500: color_o = 12'b000011110000;
		12'd501: color_o = 12'b000011110000;
		12'd502: color_o = 12'b000011110000;
		12'd503: color_o = 12'b000011110000;
		12'd504: color_o = 12'b000011110000;
		12'd505: color_o = 12'b000011110000;
		12'd506: color_o = 12'b000011110000;
		12'd507: color_o = 12'b000011110000;
		12'd508: color_o = 12'b000011110000;
		12'd509: color_o = 12'b000011110000;
		12'd510: color_o = 12'b000011110000;
		12'd511: color_o = 12'b000011110000;
		12'd512: color_o = 12'b000011110000;
		12'd513: color_o = 12'b000011110000;
		12'd514: color_o = 12'b000011110000;
		12'd515: color_o = 12'b000011110000;
		12'd516: color_o = 12'b000011110000;
		12'd517: color_o = 12'b000011110000;
		12'd518: color_o = 12'b000011110000;
		12'd519: color_o = 12'b000011110000;
		12'd520: color_o = 12'b000000000000;
		12'd521: color_o = 12'b000000000000;
		12'd522: color_o = 12'b000000000000;
		12'd523: color_o = 12'b000000000000;
		12'd524: color_o = 12'b000000000000;
		12'd525: color_o = 12'b000000000000;
		12'd526: color_o = 12'b000000000000;
		12'd527: color_o = 12'b000000000000;
		12'd528: color_o = 12'b100000000001;
		12'd529: color_o = 12'b100000000001;
		12'd530: color_o = 12'b000000000000;
		12'd531: color_o = 12'b000000000000;
		12'd532: color_o = 12'b000000000000;
		12'd533: color_o = 12'b000000000000;
		12'd534: color_o = 12'b000011110000;
		12'd535: color_o = 12'b000011110000;
		12'd536: color_o = 12'b000011110000;
		12'd537: color_o = 12'b000011110000;
		12'd538: color_o = 12'b000011110000;
		12'd539: color_o = 12'b000011110000;
		12'd540: color_o = 12'b000011110000;
		12'd541: color_o = 12'b000011110000;
		12'd542: color_o = 12'b000011110000;
		12'd543: color_o = 12'b000011110000;
		12'd544: color_o = 12'b000011110000;
		12'd545: color_o = 12'b000011110000;
		12'd546: color_o = 12'b000011110000;
		12'd547: color_o = 12'b000011110000;
		12'd548: color_o = 12'b000011110000;
		12'd549: color_o = 12'b000011110000;
		12'd550: color_o = 12'b000011110000;
		12'd551: color_o = 12'b000011110000;
		12'd552: color_o = 12'b000000000000;
		12'd553: color_o = 12'b100000000001;
		12'd554: color_o = 12'b100000000001;
		12'd555: color_o = 12'b100000000001;
		12'd556: color_o = 12'b000000000000;
		12'd557: color_o = 12'b100000000001;
		12'd558: color_o = 12'b100000000001;
		12'd559: color_o = 12'b100000000001;
		12'd560: color_o = 12'b100000000001;
		12'd561: color_o = 12'b000000000000;
		12'd562: color_o = 12'b000000000000;
		12'd563: color_o = 12'b100000000001;
		12'd564: color_o = 12'b100000000001;
		12'd565: color_o = 12'b000000000000;
		12'd566: color_o = 12'b000000000000;
		12'd567: color_o = 12'b000011110000;
		12'd568: color_o = 12'b000011110000;
		12'd569: color_o = 12'b000011110000;
		12'd570: color_o = 12'b000011110000;
		12'd571: color_o = 12'b000011110000;
		12'd572: color_o = 12'b000011110000;
		12'd573: color_o = 12'b000011110000;
		12'd574: color_o = 12'b000011110000;
		12'd575: color_o = 12'b000011110000;
		12'd576: color_o = 12'b000011110000;
		12'd577: color_o = 12'b000011110000;
		12'd578: color_o = 12'b000011110000;
		12'd579: color_o = 12'b000011110000;
		12'd580: color_o = 12'b000011110000;
		12'd581: color_o = 12'b000011110000;
		12'd582: color_o = 12'b000011110000;
		12'd583: color_o = 12'b000011110000;
		12'd584: color_o = 12'b000000000000;
		12'd585: color_o = 12'b100000000001;
		12'd586: color_o = 12'b100000000001;
		12'd587: color_o = 12'b100000000001;
		12'd588: color_o = 12'b000000000000;
		12'd589: color_o = 12'b100000000001;
		12'd590: color_o = 12'b100000000001;
		12'd591: color_o = 12'b100000000001;
		12'd592: color_o = 12'b000000000000;
		12'd593: color_o = 12'b000000000000;
		12'd594: color_o = 12'b100000000001;
		12'd595: color_o = 12'b100000000001;
		12'd596: color_o = 12'b100000000001;
		12'd597: color_o = 12'b100000000001;
		12'd598: color_o = 12'b000000000000;
		12'd599: color_o = 12'b000000000000;
		12'd600: color_o = 12'b000011110000;
		12'd601: color_o = 12'b000011110000;
		12'd602: color_o = 12'b000011110000;
		12'd603: color_o = 12'b000011110000;
		12'd604: color_o = 12'b000011110000;
		12'd605: color_o = 12'b000011110000;
		12'd606: color_o = 12'b000011110000;
		12'd607: color_o = 12'b000011110000;
		12'd608: color_o = 12'b000011110000;
		12'd609: color_o = 12'b000011110000;
		12'd610: color_o = 12'b000011110000;
		12'd611: color_o = 12'b000011110000;
		12'd612: color_o = 12'b000011110000;
		12'd613: color_o = 12'b000011110000;
		12'd614: color_o = 12'b000011110000;
		12'd615: color_o = 12'b000000000000;
		12'd616: color_o = 12'b000000000000;
		12'd617: color_o = 12'b100000000001;
		12'd618: color_o = 12'b100000000001;
		12'd619: color_o = 12'b000000000000;
		12'd620: color_o = 12'b000000000000;
		12'd621: color_o = 12'b000000000000;
		12'd622: color_o = 12'b100000000001;
		12'd623: color_o = 12'b000000000000;
		12'd624: color_o = 12'b000000000000;
		12'd625: color_o = 12'b100000000001;
		12'd626: color_o = 12'b100000000001;
		12'd627: color_o = 12'b100000000001;
		12'd628: color_o = 12'b100000000001;
		12'd629: color_o = 12'b100000000001;
		12'd630: color_o = 12'b000000000000;
		12'd631: color_o = 12'b000000000000;
		12'd632: color_o = 12'b000011110000;
		12'd633: color_o = 12'b000011110000;
		12'd634: color_o = 12'b000011110000;
		12'd635: color_o = 12'b000011110000;
		12'd636: color_o = 12'b000011110000;
		12'd637: color_o = 12'b000011110000;
		12'd638: color_o = 12'b000011110000;
		12'd639: color_o = 12'b000011110000;
		12'd640: color_o = 12'b000011110000;
		12'd641: color_o = 12'b000011110000;
		12'd642: color_o = 12'b000011110000;
		12'd643: color_o = 12'b000011110000;
		12'd644: color_o = 12'b000011110000;
		12'd645: color_o = 12'b000011110000;
		12'd646: color_o = 12'b000000000000;
		12'd647: color_o = 12'b000000000000;
		12'd648: color_o = 12'b100000000001;
		12'd649: color_o = 12'b000000000000;
		12'd650: color_o = 12'b100000000001;
		12'd651: color_o = 12'b100000000001;
		12'd652: color_o = 12'b000000000000;
		12'd653: color_o = 12'b000000000000;
		12'd654: color_o = 12'b100000000001;
		12'd655: color_o = 12'b000000000000;
		12'd656: color_o = 12'b100000000001;
		12'd657: color_o = 12'b100000000001;
		12'd658: color_o = 12'b100000000001;
		12'd659: color_o = 12'b100000000001;
		12'd660: color_o = 12'b100000000001;
		12'd661: color_o = 12'b100000000001;
		12'd662: color_o = 12'b000000000000;
		12'd663: color_o = 12'b000000000000;
		12'd664: color_o = 12'b000011110000;
		12'd665: color_o = 12'b000011110000;
		12'd666: color_o = 12'b000011110000;
		12'd667: color_o = 12'b000011110000;
		12'd668: color_o = 12'b000011110000;
		12'd669: color_o = 12'b000011110000;
		12'd670: color_o = 12'b000011110000;
		12'd671: color_o = 12'b000011110000;
		12'd672: color_o = 12'b000011110000;
		12'd673: color_o = 12'b000011110000;
		12'd674: color_o = 12'b000011110000;
		12'd675: color_o = 12'b000011110000;
		12'd676: color_o = 12'b000011110000;
		12'd677: color_o = 12'b000011110000;
		12'd678: color_o = 12'b000000000000;
		12'd679: color_o = 12'b000000000000;
		12'd680: color_o = 12'b000000000000;
		12'd681: color_o = 12'b000000000000;
		12'd682: color_o = 12'b000000000000;
		12'd683: color_o = 12'b000000000000;
		12'd684: color_o = 12'b000000000000;
		12'd685: color_o = 12'b000000000000;
		12'd686: color_o = 12'b000000000000;
		12'd687: color_o = 12'b000000000000;
		12'd688: color_o = 12'b000000000000;
		12'd689: color_o = 12'b000000000000;
		12'd690: color_o = 12'b000000000000;
		12'd691: color_o = 12'b000000000000;
		12'd692: color_o = 12'b000000000000;
		12'd693: color_o = 12'b000000000000;
		12'd694: color_o = 12'b000000000000;
		12'd695: color_o = 12'b000000000000;
		12'd696: color_o = 12'b000011110000;
		12'd697: color_o = 12'b000011110000;
		12'd698: color_o = 12'b000011110000;
		12'd699: color_o = 12'b000011110000;
		12'd700: color_o = 12'b000011110000;
		12'd701: color_o = 12'b000011110000;
		12'd702: color_o = 12'b000011110000;
		12'd703: color_o = 12'b000011110000;
		12'd704: color_o = 12'b000011110000;
		12'd705: color_o = 12'b000011110000;
		12'd706: color_o = 12'b000011110000;
		12'd707: color_o = 12'b000011110000;
		12'd708: color_o = 12'b000011110000;
		12'd709: color_o = 12'b000011110000;
		12'd710: color_o = 12'b000011110000;
		12'd711: color_o = 12'b000011110000;
		12'd712: color_o = 12'b000011110000;
		12'd713: color_o = 12'b000011110000;
		12'd714: color_o = 12'b000011110000;
		12'd715: color_o = 12'b000011110000;
		12'd716: color_o = 12'b000000000000;
		12'd717: color_o = 12'b000000000000;
		12'd718: color_o = 12'b000000000000;
		12'd719: color_o = 12'b000000000000;
		12'd720: color_o = 12'b000011110000;
		12'd721: color_o = 12'b000011110000;
		12'd722: color_o = 12'b000011110000;
		12'd723: color_o = 12'b000011110000;
		12'd724: color_o = 12'b000011110000;
		12'd725: color_o = 12'b000011110000;
		12'd726: color_o = 12'b000011110000;
		12'd727: color_o = 12'b000011110000;
		12'd728: color_o = 12'b000011110000;
		12'd729: color_o = 12'b000011110000;
		12'd730: color_o = 12'b000011110000;
		12'd731: color_o = 12'b000011110000;
		12'd732: color_o = 12'b000011110000;
		12'd733: color_o = 12'b000011110000;
		12'd734: color_o = 12'b000011110000;
		12'd735: color_o = 12'b000011110000;
		12'd736: color_o = 12'b000011110000;
		12'd737: color_o = 12'b000011110000;
		12'd738: color_o = 12'b000011110000;
		12'd739: color_o = 12'b000011110000;
		12'd740: color_o = 12'b000011110000;
		12'd741: color_o = 12'b000011110000;
		12'd742: color_o = 12'b000011110000;
		12'd743: color_o = 12'b000011110000;
		12'd744: color_o = 12'b000011110000;
		12'd745: color_o = 12'b000011110000;
		12'd746: color_o = 12'b000011110000;
		12'd747: color_o = 12'b000011110000;
		12'd748: color_o = 12'b000011110000;
		12'd749: color_o = 12'b000011110000;
		12'd750: color_o = 12'b000011110000;
		12'd751: color_o = 12'b000011110000;
		12'd752: color_o = 12'b000011110000;
		12'd753: color_o = 12'b000011110000;
		12'd754: color_o = 12'b000011110000;
		12'd755: color_o = 12'b000011110000;
		12'd756: color_o = 12'b000011110000;
		12'd757: color_o = 12'b000011110000;
		12'd758: color_o = 12'b000011110000;
		12'd759: color_o = 12'b000011110000;
		12'd760: color_o = 12'b000011110000;
		12'd761: color_o = 12'b000011110000;
		12'd762: color_o = 12'b000011110000;
		12'd763: color_o = 12'b000011110000;
		12'd764: color_o = 12'b000011110000;
		12'd765: color_o = 12'b000011110000;
		12'd766: color_o = 12'b000011110000;
		12'd767: color_o = 12'b000011110000;
		12'd768: color_o = 12'b000011110000;
		12'd769: color_o = 12'b000000000000;
		12'd770: color_o = 12'b000000000000;
		12'd771: color_o = 12'b000000000000;
		12'd772: color_o = 12'b000000000000;
		12'd773: color_o = 12'b100000000001;
		12'd774: color_o = 12'b100000000001;
		12'd775: color_o = 12'b100000000000;
		12'd776: color_o = 12'b100000000000;
		12'd777: color_o = 12'b100000000000;
		12'd778: color_o = 12'b000000000000;
		12'd779: color_o = 12'b000000000000;
		12'd780: color_o = 12'b000000000000;
		12'd781: color_o = 12'b000000000000;
		12'd782: color_o = 12'b000000000000;
		12'd783: color_o = 12'b000000000000;
		12'd784: color_o = 12'b000000000000;
		12'd785: color_o = 12'b000000000000;
		12'd786: color_o = 12'b100000000000;
		12'd787: color_o = 12'b100000000000;
		12'd788: color_o = 12'b100000000000;
		12'd789: color_o = 12'b100000000001;
		12'd790: color_o = 12'b000000000000;
		12'd791: color_o = 12'b000011110000;
		12'd792: color_o = 12'b000011110000;
		12'd793: color_o = 12'b000011110000;
		12'd794: color_o = 12'b000011110000;
		12'd795: color_o = 12'b000011110000;
		12'd796: color_o = 12'b000011110000;
		12'd797: color_o = 12'b000011110000;
		12'd798: color_o = 12'b000011110000;
		12'd799: color_o = 12'b000011110000;
		12'd800: color_o = 12'b000011110000;
		12'd801: color_o = 12'b000000000000;
		12'd802: color_o = 12'b000000000000;
		12'd803: color_o = 12'b000000000000;
		12'd804: color_o = 12'b000000000000;
		12'd805: color_o = 12'b100000000001;
		12'd806: color_o = 12'b100000000001;
		12'd807: color_o = 12'b100000000001;
		12'd808: color_o = 12'b100000000001;
		12'd809: color_o = 12'b000000000000;
		12'd810: color_o = 12'b000000000000;
		12'd811: color_o = 12'b000000000000;
		12'd812: color_o = 12'b000000000000;
		12'd813: color_o = 12'b000000000000;
		12'd814: color_o = 12'b100000000000;
		12'd815: color_o = 12'b100000000000;
		12'd816: color_o = 12'b100000000000;
		12'd817: color_o = 12'b100000000000;
		12'd818: color_o = 12'b000000000000;
		12'd819: color_o = 12'b100000000000;
		12'd820: color_o = 12'b100000000001;
		12'd821: color_o = 12'b100000000001;
		12'd822: color_o = 12'b000000000000;
		12'd823: color_o = 12'b000011110000;
		12'd824: color_o = 12'b000011110000;
		12'd825: color_o = 12'b000011110000;
		12'd826: color_o = 12'b000011110000;
		12'd827: color_o = 12'b000011110000;
		12'd828: color_o = 12'b000011110000;
		12'd829: color_o = 12'b000011110000;
		12'd830: color_o = 12'b000011110000;
		12'd831: color_o = 12'b000011110000;
		12'd832: color_o = 12'b000011110000;
		12'd833: color_o = 12'b000000000000;
		12'd834: color_o = 12'b000000000000;
		12'd835: color_o = 12'b000000000000;
		12'd836: color_o = 12'b000000000000;
		12'd837: color_o = 12'b000000000000;
		12'd838: color_o = 12'b000000000000;
		12'd839: color_o = 12'b100000000000;
		12'd840: color_o = 12'b100000000001;
		12'd841: color_o = 12'b100000000001;
		12'd842: color_o = 12'b100000000000;
		12'd843: color_o = 12'b100000000000;
		12'd844: color_o = 12'b100000000000;
		12'd845: color_o = 12'b100000000000;
		12'd846: color_o = 12'b010000000000;
		12'd847: color_o = 12'b010000000000;
		12'd848: color_o = 12'b010000000000;
		12'd849: color_o = 12'b010000000000;
		12'd850: color_o = 12'b000000000000;
		12'd851: color_o = 12'b000000000000;
		12'd852: color_o = 12'b000000000000;
		12'd853: color_o = 12'b000000000000;
		12'd854: color_o = 12'b000000000000;
		12'd855: color_o = 12'b000011110000;
		12'd856: color_o = 12'b000011110000;
		12'd857: color_o = 12'b000011110000;
		12'd858: color_o = 12'b000011110000;
		12'd859: color_o = 12'b000011110000;
		12'd860: color_o = 12'b000011110000;
		12'd861: color_o = 12'b000011110000;
		12'd862: color_o = 12'b000011110000;
		12'd863: color_o = 12'b000011110000;
		12'd864: color_o = 12'b000011110000;
		12'd865: color_o = 12'b000011110000;
		12'd866: color_o = 12'b000000000000;
		12'd867: color_o = 12'b000000000000;
		12'd868: color_o = 12'b100000000001;
		12'd869: color_o = 12'b100000000001;
		12'd870: color_o = 12'b000000000000;
		12'd871: color_o = 12'b000000000000;
		12'd872: color_o = 12'b000000000000;
		12'd873: color_o = 12'b000000000000;
		12'd874: color_o = 12'b100000000000;
		12'd875: color_o = 12'b010000000000;
		12'd876: color_o = 12'b010000000000;
		12'd877: color_o = 12'b010000000000;
		12'd878: color_o = 12'b010000000000;
		12'd879: color_o = 12'b010000000000;
		12'd880: color_o = 12'b000000000000;
		12'd881: color_o = 12'b000000000000;
		12'd882: color_o = 12'b000000000000;
		12'd883: color_o = 12'b010000000000;
		12'd884: color_o = 12'b010000000000;
		12'd885: color_o = 12'b000000000000;
		12'd886: color_o = 12'b000011110000;
		12'd887: color_o = 12'b000011110000;
		12'd888: color_o = 12'b000011110000;
		12'd889: color_o = 12'b000011110000;
		12'd890: color_o = 12'b000011110000;
		12'd891: color_o = 12'b000011110000;
		12'd892: color_o = 12'b000011110000;
		12'd893: color_o = 12'b000011110000;
		12'd894: color_o = 12'b000011110000;
		12'd895: color_o = 12'b000011110000;
		12'd896: color_o = 12'b000011110000;
		12'd897: color_o = 12'b000011110000;
		12'd898: color_o = 12'b000000000000;
		12'd899: color_o = 12'b100000000001;
		12'd900: color_o = 12'b100000000001;
		12'd901: color_o = 12'b000000000000;
		12'd902: color_o = 12'b000000000000;
		12'd903: color_o = 12'b000000000000;
		12'd904: color_o = 12'b000000000000;
		12'd905: color_o = 12'b000000000000;
		12'd906: color_o = 12'b000000000000;
		12'd907: color_o = 12'b000000000000;
		12'd908: color_o = 12'b000000000000;
		12'd909: color_o = 12'b000000000000;
		12'd910: color_o = 12'b000000000000;
		12'd911: color_o = 12'b000000000000;
		12'd912: color_o = 12'b000000000000;
		12'd913: color_o = 12'b000000000000;
		12'd914: color_o = 12'b100000000001;
		12'd915: color_o = 12'b100000000001;
		12'd916: color_o = 12'b000000000000;
		12'd917: color_o = 12'b000000000000;
		12'd918: color_o = 12'b000011110000;
		12'd919: color_o = 12'b000011110000;
		12'd920: color_o = 12'b000011110000;
		12'd921: color_o = 12'b000011110000;
		12'd922: color_o = 12'b000011110000;
		12'd923: color_o = 12'b000011110000;
		12'd924: color_o = 12'b000011110000;
		12'd925: color_o = 12'b000011110000;
		12'd926: color_o = 12'b000011110000;
		12'd927: color_o = 12'b000011110000;
		12'd928: color_o = 12'b000011110000;
		12'd929: color_o = 12'b000011110000;
		12'd930: color_o = 12'b000000000000;
		12'd931: color_o = 12'b000000000000;
		12'd932: color_o = 12'b100000000001;
		12'd933: color_o = 12'b100000000001;
		12'd934: color_o = 12'b100000000001;
		12'd935: color_o = 12'b100000000001;
		12'd936: color_o = 12'b100000000001;
		12'd937: color_o = 12'b100000000001;
		12'd938: color_o = 12'b100000000001;
		12'd939: color_o = 12'b100000000001;
		12'd940: color_o = 12'b100000000001;
		12'd941: color_o = 12'b100000000001;
		12'd942: color_o = 12'b100000000001;
		12'd943: color_o = 12'b100000000001;
		12'd944: color_o = 12'b100000000001;
		12'd945: color_o = 12'b100000000001;
		12'd946: color_o = 12'b100000000001;
		12'd947: color_o = 12'b100000000001;
		12'd948: color_o = 12'b100000000001;
		12'd949: color_o = 12'b100000000001;
		12'd950: color_o = 12'b000000000000;
		12'd951: color_o = 12'b000011110000;
		12'd952: color_o = 12'b000011110000;
		12'd953: color_o = 12'b000011110000;
		12'd954: color_o = 12'b000011110000;
		12'd955: color_o = 12'b000011110000;
		12'd956: color_o = 12'b000011110000;
		12'd957: color_o = 12'b000011110000;
		12'd958: color_o = 12'b000011110000;
		12'd959: color_o = 12'b000011110000;
		12'd960: color_o = 12'b000011110000;
		12'd961: color_o = 12'b000011110000;
		12'd962: color_o = 12'b000000000000;
		12'd963: color_o = 12'b000000000000;
		12'd964: color_o = 12'b100000000001;
		12'd965: color_o = 12'b100000000001;
		12'd966: color_o = 12'b100000000001;
		12'd967: color_o = 12'b000000000000;
		12'd968: color_o = 12'b000000000000;
		12'd969: color_o = 12'b100000000001;
		12'd970: color_o = 12'b100000000001;
		12'd971: color_o = 12'b100000000001;
		12'd972: color_o = 12'b100000000001;
		12'd973: color_o = 12'b100000000001;
		12'd974: color_o = 12'b100000000001;
		12'd975: color_o = 12'b100000000001;
		12'd976: color_o = 12'b100000000001;
		12'd977: color_o = 12'b100000000001;
		12'd978: color_o = 12'b100000000001;
		12'd979: color_o = 12'b100000000001;
		12'd980: color_o = 12'b000000000000;
		12'd981: color_o = 12'b000000000000;
		12'd982: color_o = 12'b000000000000;
		12'd983: color_o = 12'b000000000000;
		12'd984: color_o = 12'b000011110000;
		12'd985: color_o = 12'b000011110000;
		12'd986: color_o = 12'b000011110000;
		12'd987: color_o = 12'b000011110000;
		12'd988: color_o = 12'b000011110000;
		12'd989: color_o = 12'b000011110000;
		12'd990: color_o = 12'b000011110000;
		12'd991: color_o = 12'b000011110000;
		12'd992: color_o = 12'b000011110000;
		12'd993: color_o = 12'b000011110000;
		12'd994: color_o = 12'b000000000000;
		12'd995: color_o = 12'b000000000000;
		12'd996: color_o = 12'b000000000000;
		12'd997: color_o = 12'b100000000001;
		12'd998: color_o = 12'b100000000001;
		12'd999: color_o = 12'b010000000000;
		12'd1000: color_o = 12'b000000000000;
		12'd1001: color_o = 12'b100000000001;
		12'd1002: color_o = 12'b000000000000;
		12'd1003: color_o = 12'b000000000000;
		12'd1004: color_o = 12'b100000000001;
		12'd1005: color_o = 12'b100000000001;
		12'd1006: color_o = 12'b100000000001;
		12'd1007: color_o = 12'b100000000001;
		12'd1008: color_o = 12'b100000000001;
		12'd1009: color_o = 12'b100000000001;
		12'd1010: color_o = 12'b000000000000;
		12'd1011: color_o = 12'b000000000000;
		12'd1012: color_o = 12'b000000000000;
		12'd1013: color_o = 12'b100000000001;
		12'd1014: color_o = 12'b100000000001;
		12'd1015: color_o = 12'b000000000000;
		12'd1016: color_o = 12'b000011110000;
		12'd1017: color_o = 12'b000011110000;
		12'd1018: color_o = 12'b000011110000;
		12'd1019: color_o = 12'b000011110000;
		12'd1020: color_o = 12'b000011110000;
		12'd1021: color_o = 12'b000011110000;
		12'd1022: color_o = 12'b000011110000;
		12'd1023: color_o = 12'b000011110000;
		12'd1024: color_o = 12'b000011110000;
		12'd1025: color_o = 12'b000011110000;
		12'd1026: color_o = 12'b000011110000;
		12'd1027: color_o = 12'b000000000000;
		12'd1028: color_o = 12'b000000000000;
		12'd1029: color_o = 12'b000000000000;
		12'd1030: color_o = 12'b000000000000;
		12'd1031: color_o = 12'b000000000000;
		12'd1032: color_o = 12'b000000000000;
		12'd1033: color_o = 12'b100000000001;
		12'd1034: color_o = 12'b010000000000;
		12'd1035: color_o = 12'b000000000000;
		12'd1036: color_o = 12'b100000000001;
		12'd1037: color_o = 12'b100000000001;
		12'd1038: color_o = 12'b100000000001;
		12'd1039: color_o = 12'b100000000001;
		12'd1040: color_o = 12'b100000000001;
		12'd1041: color_o = 12'b100000000001;
		12'd1042: color_o = 12'b100000000001;
		12'd1043: color_o = 12'b100000000001;
		12'd1044: color_o = 12'b100000000001;
		12'd1045: color_o = 12'b100000000001;
		12'd1046: color_o = 12'b100000000001;
		12'd1047: color_o = 12'b100000000001;
		12'd1048: color_o = 12'b000000000000;
		12'd1049: color_o = 12'b000011110000;
		12'd1050: color_o = 12'b000011110000;
		12'd1051: color_o = 12'b000011110000;
		12'd1052: color_o = 12'b000011110000;
		12'd1053: color_o = 12'b000011110000;
		12'd1054: color_o = 12'b000011110000;
		12'd1055: color_o = 12'b000011110000;
		12'd1056: color_o = 12'b000011110000;
		12'd1057: color_o = 12'b000011110000;
		12'd1058: color_o = 12'b000011110000;
		12'd1059: color_o = 12'b000000000000;
		12'd1060: color_o = 12'b000000000000;
		12'd1061: color_o = 12'b000000000000;
		12'd1062: color_o = 12'b000000000000;
		12'd1063: color_o = 12'b000000000000;
		12'd1064: color_o = 12'b000000000000;
		12'd1065: color_o = 12'b100000000001;
		12'd1066: color_o = 12'b010000000000;
		12'd1067: color_o = 12'b000000000000;
		12'd1068: color_o = 12'b100000000001;
		12'd1069: color_o = 12'b100000000001;
		12'd1070: color_o = 12'b100000000001;
		12'd1071: color_o = 12'b100000000001;
		12'd1072: color_o = 12'b100000000001;
		12'd1073: color_o = 12'b100000000001;
		12'd1074: color_o = 12'b000000000000;
		12'd1075: color_o = 12'b100000000001;
		12'd1076: color_o = 12'b100000000001;
		12'd1077: color_o = 12'b100000000001;
		12'd1078: color_o = 12'b100000000001;
		12'd1079: color_o = 12'b100000000001;
		12'd1080: color_o = 12'b000000000000;
		12'd1081: color_o = 12'b000011110000;
		12'd1082: color_o = 12'b000011110000;
		12'd1083: color_o = 12'b000011110000;
		12'd1084: color_o = 12'b000011110000;
		12'd1085: color_o = 12'b000011110000;
		12'd1086: color_o = 12'b000011110000;
		12'd1087: color_o = 12'b000011110000;
		12'd1088: color_o = 12'b000011110000;
		12'd1089: color_o = 12'b000011110000;
		12'd1090: color_o = 12'b000011110000;
		12'd1091: color_o = 12'b000000000000;
		12'd1092: color_o = 12'b000000000000;
		12'd1093: color_o = 12'b000000000000;
		12'd1094: color_o = 12'b000000000000;
		12'd1095: color_o = 12'b010000000000;
		12'd1096: color_o = 12'b000000000000;
		12'd1097: color_o = 12'b000000000000;
		12'd1098: color_o = 12'b000000000000;
		12'd1099: color_o = 12'b000000000000;
		12'd1100: color_o = 12'b000000000000;
		12'd1101: color_o = 12'b100000000001;
		12'd1102: color_o = 12'b100000000001;
		12'd1103: color_o = 12'b100000000001;
		12'd1104: color_o = 12'b100000000001;
		12'd1105: color_o = 12'b100000000001;
		12'd1106: color_o = 12'b000000000000;
		12'd1107: color_o = 12'b100000000001;
		12'd1108: color_o = 12'b100000000001;
		12'd1109: color_o = 12'b100000000001;
		12'd1110: color_o = 12'b100000000001;
		12'd1111: color_o = 12'b100000000001;
		12'd1112: color_o = 12'b000000000000;
		12'd1113: color_o = 12'b000011110000;
		12'd1114: color_o = 12'b000011110000;
		12'd1115: color_o = 12'b000011110000;
		12'd1116: color_o = 12'b000011110000;
		12'd1117: color_o = 12'b000011110000;
		12'd1118: color_o = 12'b000011110000;
		12'd1119: color_o = 12'b000011110000;
		12'd1120: color_o = 12'b000011110000;
		12'd1121: color_o = 12'b000011110000;
		12'd1122: color_o = 12'b000000000000;
		12'd1123: color_o = 12'b000000000000;
		12'd1124: color_o = 12'b000000000000;
		12'd1125: color_o = 12'b000000000000;
		12'd1126: color_o = 12'b000000000000;
		12'd1127: color_o = 12'b010000000000;
		12'd1128: color_o = 12'b010000000000;
		12'd1129: color_o = 12'b000000000000;
		12'd1130: color_o = 12'b000000000000;
		12'd1131: color_o = 12'b000000000000;
		12'd1132: color_o = 12'b000000000000;
		12'd1133: color_o = 12'b100000000001;
		12'd1134: color_o = 12'b100000000001;
		12'd1135: color_o = 12'b100000000001;
		12'd1136: color_o = 12'b100000000001;
		12'd1137: color_o = 12'b100000000001;
		12'd1138: color_o = 12'b000000000000;
		12'd1139: color_o = 12'b010000000000;
		12'd1140: color_o = 12'b010000000000;
		12'd1141: color_o = 12'b100000000001;
		12'd1142: color_o = 12'b010000000000;
		12'd1143: color_o = 12'b000000000000;
		12'd1144: color_o = 12'b000000000000;
		12'd1145: color_o = 12'b000011110000;
		12'd1146: color_o = 12'b000011110000;
		12'd1147: color_o = 12'b000011110000;
		12'd1148: color_o = 12'b000011110000;
		12'd1149: color_o = 12'b000011110000;
		12'd1150: color_o = 12'b000011110000;
		12'd1151: color_o = 12'b000011110000;
		12'd1152: color_o = 12'b000011110000;
		12'd1153: color_o = 12'b000011110000;
		12'd1154: color_o = 12'b000000000000;
		12'd1155: color_o = 12'b000000000000;
		12'd1156: color_o = 12'b000000000000;
		12'd1157: color_o = 12'b000000000000;
		12'd1158: color_o = 12'b000000000000;
		12'd1159: color_o = 12'b000000000000;
		12'd1160: color_o = 12'b010000000000;
		12'd1161: color_o = 12'b010000000000;
		12'd1162: color_o = 12'b000000000000;
		12'd1163: color_o = 12'b000000000000;
		12'd1164: color_o = 12'b000000000000;
		12'd1165: color_o = 12'b100000000001;
		12'd1166: color_o = 12'b000000000000;
		12'd1167: color_o = 12'b000000000000;
		12'd1168: color_o = 12'b000000000000;
		12'd1169: color_o = 12'b100000000001;
		12'd1170: color_o = 12'b000000000000;
		12'd1171: color_o = 12'b000000000000;
		12'd1172: color_o = 12'b010000000000;
		12'd1173: color_o = 12'b010000000000;
		12'd1174: color_o = 12'b010000000000;
		12'd1175: color_o = 12'b000000000000;
		12'd1176: color_o = 12'b000011110000;
		12'd1177: color_o = 12'b000011110000;
		12'd1178: color_o = 12'b000011110000;
		12'd1179: color_o = 12'b000011110000;
		12'd1180: color_o = 12'b000011110000;
		12'd1181: color_o = 12'b000011110000;
		12'd1182: color_o = 12'b000011110000;
		12'd1183: color_o = 12'b000011110000;
		12'd1184: color_o = 12'b000011110000;
		12'd1185: color_o = 12'b000011110000;
		12'd1186: color_o = 12'b000000000000;
		12'd1187: color_o = 12'b000000000000;
		12'd1188: color_o = 12'b000000000000;
		12'd1189: color_o = 12'b000000000000;
		12'd1190: color_o = 12'b000000000000;
		12'd1191: color_o = 12'b000000000000;
		12'd1192: color_o = 12'b000000000000;
		12'd1193: color_o = 12'b000000000000;
		12'd1194: color_o = 12'b000000000000;
		12'd1195: color_o = 12'b000000000000;
		12'd1196: color_o = 12'b000011110000;
		12'd1197: color_o = 12'b000000000000;
		12'd1198: color_o = 12'b000000000000;
		12'd1199: color_o = 12'b000000000000;
		12'd1200: color_o = 12'b100000000001;
		12'd1201: color_o = 12'b100000000001;
		12'd1202: color_o = 12'b100000000001;
		12'd1203: color_o = 12'b100000000001;
		12'd1204: color_o = 12'b000000000000;
		12'd1205: color_o = 12'b000000000000;
		12'd1206: color_o = 12'b000000000000;
		12'd1207: color_o = 12'b000000000000;
		12'd1208: color_o = 12'b000011110000;
		12'd1209: color_o = 12'b000011110000;
		12'd1210: color_o = 12'b000011110000;
		12'd1211: color_o = 12'b000011110000;
		12'd1212: color_o = 12'b000011110000;
		12'd1213: color_o = 12'b000011110000;
		12'd1214: color_o = 12'b000011110000;
		12'd1215: color_o = 12'b000011110000;
		12'd1216: color_o = 12'b000011110000;
		12'd1217: color_o = 12'b000011110000;
		12'd1218: color_o = 12'b000000000000;
		12'd1219: color_o = 12'b000000000000;
		12'd1220: color_o = 12'b000000000000;
		12'd1221: color_o = 12'b000000000000;
		12'd1222: color_o = 12'b000000000000;
		12'd1223: color_o = 12'b000000000000;
		12'd1224: color_o = 12'b000000000000;
		12'd1225: color_o = 12'b010000000000;
		12'd1226: color_o = 12'b000000000000;
		12'd1227: color_o = 12'b000011110000;
		12'd1228: color_o = 12'b000011110000;
		12'd1229: color_o = 12'b000011110000;
		12'd1230: color_o = 12'b000000000000;
		12'd1231: color_o = 12'b000000000000;
		12'd1232: color_o = 12'b100000000001;
		12'd1233: color_o = 12'b100000000001;
		12'd1234: color_o = 12'b100000000001;
		12'd1235: color_o = 12'b100000000001;
		12'd1236: color_o = 12'b100000000001;
		12'd1237: color_o = 12'b100000000001;
		12'd1238: color_o = 12'b000000000000;
		12'd1239: color_o = 12'b000000000000;
		12'd1240: color_o = 12'b000000000000;
		12'd1241: color_o = 12'b000000000000;
		12'd1242: color_o = 12'b000011110000;
		12'd1243: color_o = 12'b000011110000;
		12'd1244: color_o = 12'b000011110000;
		12'd1245: color_o = 12'b000011110000;
		12'd1246: color_o = 12'b000011110000;
		12'd1247: color_o = 12'b000011110000;
		12'd1248: color_o = 12'b000011110000;
		12'd1249: color_o = 12'b000000000000;
		12'd1250: color_o = 12'b000000000000;
		12'd1251: color_o = 12'b000000000000;
		12'd1252: color_o = 12'b000000000000;
		12'd1253: color_o = 12'b000000000000;
		12'd1254: color_o = 12'b000000000000;
		12'd1255: color_o = 12'b000000000000;
		12'd1256: color_o = 12'b000000000000;
		12'd1257: color_o = 12'b010000000000;
		12'd1258: color_o = 12'b000011110000;
		12'd1259: color_o = 12'b000011110000;
		12'd1260: color_o = 12'b000011110000;
		12'd1261: color_o = 12'b000011110000;
		12'd1262: color_o = 12'b000011110000;
		12'd1263: color_o = 12'b000000000000;
		12'd1264: color_o = 12'b000000000000;
		12'd1265: color_o = 12'b000000000000;
		12'd1266: color_o = 12'b100000000001;
		12'd1267: color_o = 12'b100000000001;
		12'd1268: color_o = 12'b100000000001;
		12'd1269: color_o = 12'b000000000000;
		12'd1270: color_o = 12'b000000000000;
		12'd1271: color_o = 12'b000000000000;
		12'd1272: color_o = 12'b000000000000;
		12'd1273: color_o = 12'b000000000000;
		12'd1274: color_o = 12'b000000000000;
		12'd1275: color_o = 12'b000011110000;
		12'd1276: color_o = 12'b000011110000;
		12'd1277: color_o = 12'b000011110000;
		12'd1278: color_o = 12'b000011110000;
		12'd1279: color_o = 12'b000011110000;
		12'd1280: color_o = 12'b000011110000;
		12'd1281: color_o = 12'b000000000000;
		12'd1282: color_o = 12'b000000000000;
		12'd1283: color_o = 12'b000000000000;
		12'd1284: color_o = 12'b000000000000;
		12'd1285: color_o = 12'b000000000000;
		12'd1286: color_o = 12'b000000000000;
		12'd1287: color_o = 12'b000000000000;
		12'd1288: color_o = 12'b000000000000;
		12'd1289: color_o = 12'b010000000000;
		12'd1290: color_o = 12'b000000000000;
		12'd1291: color_o = 12'b000011110000;
		12'd1292: color_o = 12'b000011110000;
		12'd1293: color_o = 12'b000011110000;
		12'd1294: color_o = 12'b000011110000;
		12'd1295: color_o = 12'b000000000000;
		12'd1296: color_o = 12'b000000000000;
		12'd1297: color_o = 12'b000000000000;
		12'd1298: color_o = 12'b000000000000;
		12'd1299: color_o = 12'b000000000000;
		12'd1300: color_o = 12'b000000000000;
		12'd1301: color_o = 12'b000000000000;
		12'd1302: color_o = 12'b000000000000;
		12'd1303: color_o = 12'b100000000001;
		12'd1304: color_o = 12'b100000000001;
		12'd1305: color_o = 12'b000000000000;
		12'd1306: color_o = 12'b000000000000;
		12'd1307: color_o = 12'b000000000000;
		12'd1308: color_o = 12'b000000000000;
		12'd1309: color_o = 12'b000011110000;
		12'd1310: color_o = 12'b000011110000;
		12'd1311: color_o = 12'b000011110000;
		12'd1312: color_o = 12'b000000000000;
		12'd1313: color_o = 12'b000000000000;
		12'd1314: color_o = 12'b000000000000;
		12'd1315: color_o = 12'b000000000000;
		12'd1316: color_o = 12'b000000000000;
		12'd1317: color_o = 12'b000000000000;
		12'd1318: color_o = 12'b100000000001;
		12'd1319: color_o = 12'b100000000001;
		12'd1320: color_o = 12'b100000000001;
		12'd1321: color_o = 12'b100000000001;
		12'd1322: color_o = 12'b000000000000;
		12'd1323: color_o = 12'b000000000000;
		12'd1324: color_o = 12'b000011110000;
		12'd1325: color_o = 12'b000011110000;
		12'd1326: color_o = 12'b000011110000;
		12'd1327: color_o = 12'b000000000000;
		12'd1328: color_o = 12'b100000000001;
		12'd1329: color_o = 12'b100000000001;
		12'd1330: color_o = 12'b100000000001;
		12'd1331: color_o = 12'b000000000000;
		12'd1332: color_o = 12'b100000000001;
		12'd1333: color_o = 12'b100000000001;
		12'd1334: color_o = 12'b100000000001;
		12'd1335: color_o = 12'b100000000001;
		12'd1336: color_o = 12'b000000000000;
		12'd1337: color_o = 12'b000000000000;
		12'd1338: color_o = 12'b100000000001;
		12'd1339: color_o = 12'b100000000001;
		12'd1340: color_o = 12'b000000000000;
		12'd1341: color_o = 12'b000000000000;
		12'd1342: color_o = 12'b000011110000;
		12'd1343: color_o = 12'b000011110000;
		12'd1344: color_o = 12'b000011110000;
		12'd1345: color_o = 12'b000000000000;
		12'd1346: color_o = 12'b000000000000;
		12'd1347: color_o = 12'b000000000000;
		12'd1348: color_o = 12'b000000000000;
		12'd1349: color_o = 12'b000000000000;
		12'd1350: color_o = 12'b000000000000;
		12'd1351: color_o = 12'b000000000000;
		12'd1352: color_o = 12'b000000000000;
		12'd1353: color_o = 12'b000000000000;
		12'd1354: color_o = 12'b000000000000;
		12'd1355: color_o = 12'b000000000000;
		12'd1356: color_o = 12'b000000000000;
		12'd1357: color_o = 12'b000011110000;
		12'd1358: color_o = 12'b000011110000;
		12'd1359: color_o = 12'b000000000000;
		12'd1360: color_o = 12'b100000000001;
		12'd1361: color_o = 12'b100000000001;
		12'd1362: color_o = 12'b100000000001;
		12'd1363: color_o = 12'b000000000000;
		12'd1364: color_o = 12'b100000000001;
		12'd1365: color_o = 12'b100000000001;
		12'd1366: color_o = 12'b100000000001;
		12'd1367: color_o = 12'b000000000000;
		12'd1368: color_o = 12'b000000000000;
		12'd1369: color_o = 12'b100000000001;
		12'd1370: color_o = 12'b100000000001;
		12'd1371: color_o = 12'b100000000001;
		12'd1372: color_o = 12'b100000000001;
		12'd1373: color_o = 12'b000000000000;
		12'd1374: color_o = 12'b000000000000;
		12'd1375: color_o = 12'b000011110000;
		12'd1376: color_o = 12'b000011110000;
		12'd1377: color_o = 12'b000011110000;
		12'd1378: color_o = 12'b000000000000;
		12'd1379: color_o = 12'b000000000000;
		12'd1380: color_o = 12'b000000000000;
		12'd1381: color_o = 12'b000000000000;
		12'd1382: color_o = 12'b000000000000;
		12'd1383: color_o = 12'b000000000000;
		12'd1384: color_o = 12'b100000000001;
		12'd1385: color_o = 12'b000000000000;
		12'd1386: color_o = 12'b000000000000;
		12'd1387: color_o = 12'b000000000000;
		12'd1388: color_o = 12'b000000000000;
		12'd1389: color_o = 12'b000011110000;
		12'd1390: color_o = 12'b000000000000;
		12'd1391: color_o = 12'b000000000000;
		12'd1392: color_o = 12'b100000000001;
		12'd1393: color_o = 12'b100000000001;
		12'd1394: color_o = 12'b000000000000;
		12'd1395: color_o = 12'b000000000000;
		12'd1396: color_o = 12'b000000000000;
		12'd1397: color_o = 12'b100000000001;
		12'd1398: color_o = 12'b000000000000;
		12'd1399: color_o = 12'b000000000000;
		12'd1400: color_o = 12'b100000000001;
		12'd1401: color_o = 12'b100000000001;
		12'd1402: color_o = 12'b100000000001;
		12'd1403: color_o = 12'b100000000001;
		12'd1404: color_o = 12'b100000000001;
		12'd1405: color_o = 12'b000000000000;
		12'd1406: color_o = 12'b000000000000;
		12'd1407: color_o = 12'b000011110000;
		12'd1408: color_o = 12'b000011110000;
		12'd1409: color_o = 12'b000011110000;
		12'd1410: color_o = 12'b000011110000;
		12'd1411: color_o = 12'b000000000000;
		12'd1412: color_o = 12'b000000000000;
		12'd1413: color_o = 12'b000000000000;
		12'd1414: color_o = 12'b000000000000;
		12'd1415: color_o = 12'b000000000000;
		12'd1416: color_o = 12'b100000000001;
		12'd1417: color_o = 12'b000000000000;
		12'd1418: color_o = 12'b000000000000;
		12'd1419: color_o = 12'b000000000000;
		12'd1420: color_o = 12'b000000000000;
		12'd1421: color_o = 12'b000000000000;
		12'd1422: color_o = 12'b000000000000;
		12'd1423: color_o = 12'b100000000001;
		12'd1424: color_o = 12'b000000000000;
		12'd1425: color_o = 12'b100000000001;
		12'd1426: color_o = 12'b100000000001;
		12'd1427: color_o = 12'b000000000000;
		12'd1428: color_o = 12'b000000000000;
		12'd1429: color_o = 12'b100000000001;
		12'd1430: color_o = 12'b000000000000;
		12'd1431: color_o = 12'b100000000001;
		12'd1432: color_o = 12'b100000000001;
		12'd1433: color_o = 12'b100000000001;
		12'd1434: color_o = 12'b100000000001;
		12'd1435: color_o = 12'b100000000001;
		12'd1436: color_o = 12'b100000000001;
		12'd1437: color_o = 12'b000000000000;
		12'd1438: color_o = 12'b000000000000;
		12'd1439: color_o = 12'b000011110000;
		12'd1440: color_o = 12'b000011110000;
		12'd1441: color_o = 12'b000011110000;
		12'd1442: color_o = 12'b000011110000;
		12'd1443: color_o = 12'b000011110000;
		12'd1444: color_o = 12'b000011110000;
		12'd1445: color_o = 12'b000011110000;
		12'd1446: color_o = 12'b000011110000;
		12'd1447: color_o = 12'b000011110000;
		12'd1448: color_o = 12'b000011110000;
		12'd1449: color_o = 12'b000011110000;
		12'd1450: color_o = 12'b000011110000;
		12'd1451: color_o = 12'b000011110000;
		12'd1452: color_o = 12'b000011110000;
		12'd1453: color_o = 12'b000000000000;
		12'd1454: color_o = 12'b000000000000;
		12'd1455: color_o = 12'b000000000000;
		12'd1456: color_o = 12'b000000000000;
		12'd1457: color_o = 12'b000000000000;
		12'd1458: color_o = 12'b000000000000;
		12'd1459: color_o = 12'b000000000000;
		12'd1460: color_o = 12'b000000000000;
		12'd1461: color_o = 12'b000000000000;
		12'd1462: color_o = 12'b000000000000;
		12'd1463: color_o = 12'b000000000000;
		12'd1464: color_o = 12'b000000000000;
		12'd1465: color_o = 12'b000000000000;
		12'd1466: color_o = 12'b000000000000;
		12'd1467: color_o = 12'b000000000000;
		12'd1468: color_o = 12'b000000000000;
		12'd1469: color_o = 12'b000000000000;
		12'd1470: color_o = 12'b000000000000;
		12'd1471: color_o = 12'b000011110000;
		12'd1472: color_o = 12'b000011110000;
		12'd1473: color_o = 12'b000011110000;
		12'd1474: color_o = 12'b000011110000;
		12'd1475: color_o = 12'b000011110000;
		12'd1476: color_o = 12'b000011110000;
		12'd1477: color_o = 12'b000011110000;
		12'd1478: color_o = 12'b000011110000;
		12'd1479: color_o = 12'b000011110000;
		12'd1480: color_o = 12'b000011110000;
		12'd1481: color_o = 12'b000011110000;
		12'd1482: color_o = 12'b000011110000;
		12'd1483: color_o = 12'b000011110000;
		12'd1484: color_o = 12'b000011110000;
		12'd1485: color_o = 12'b000011110000;
		12'd1486: color_o = 12'b000011110000;
		12'd1487: color_o = 12'b000011110000;
		12'd1488: color_o = 12'b000011110000;
		12'd1489: color_o = 12'b000011110000;
		12'd1490: color_o = 12'b000011110000;
		12'd1491: color_o = 12'b000000000000;
		12'd1492: color_o = 12'b000000000000;
		12'd1493: color_o = 12'b000000000000;
		12'd1494: color_o = 12'b000000000000;
		12'd1495: color_o = 12'b000011110000;
		12'd1496: color_o = 12'b000011110000;
		12'd1497: color_o = 12'b000011110000;
		12'd1498: color_o = 12'b000011110000;
		12'd1499: color_o = 12'b000011110000;
		12'd1500: color_o = 12'b000011110000;
		12'd1501: color_o = 12'b000011110000;
		12'd1502: color_o = 12'b000011110000;
		12'd1503: color_o = 12'b000011110000;
		12'd1504: color_o = 12'b000011110000;
		12'd1505: color_o = 12'b000011110000;
		12'd1506: color_o = 12'b000011110000;
		12'd1507: color_o = 12'b000011110000;
		12'd1508: color_o = 12'b000011110000;
		12'd1509: color_o = 12'b000011110000;
		12'd1510: color_o = 12'b000011110000;
		12'd1511: color_o = 12'b000011110000;
		12'd1512: color_o = 12'b000011110000;
		12'd1513: color_o = 12'b000011110000;
		12'd1514: color_o = 12'b000011110000;
		12'd1515: color_o = 12'b000011110000;
		12'd1516: color_o = 12'b000011110000;
		12'd1517: color_o = 12'b000011110000;
		12'd1518: color_o = 12'b000011110000;
		12'd1519: color_o = 12'b000011110000;
		12'd1520: color_o = 12'b000011110000;
		12'd1521: color_o = 12'b000011110000;
		12'd1522: color_o = 12'b000011110000;
		12'd1523: color_o = 12'b000011110000;
		12'd1524: color_o = 12'b000011110000;
		12'd1525: color_o = 12'b000011110000;
		12'd1526: color_o = 12'b000011110000;
		12'd1527: color_o = 12'b000011110000;
		12'd1528: color_o = 12'b000011110000;
		12'd1529: color_o = 12'b000011110000;
		12'd1530: color_o = 12'b000011110000;
		12'd1531: color_o = 12'b000011110000;
		12'd1532: color_o = 12'b000011110000;
		12'd1533: color_o = 12'b000011110000;
		12'd1534: color_o = 12'b000011110000;
		12'd1535: color_o = 12'b000011110000;
		12'd1536: color_o = 12'b000011110000;
		12'd1537: color_o = 12'b000011110000;
		12'd1538: color_o = 12'b000000000000;
		12'd1539: color_o = 12'b000000000000;
		12'd1540: color_o = 12'b000000000000;
		12'd1541: color_o = 12'b100000000001;
		12'd1542: color_o = 12'b100000000001;
		12'd1543: color_o = 12'b100000000000;
		12'd1544: color_o = 12'b100000000000;
		12'd1545: color_o = 12'b100000000000;
		12'd1546: color_o = 12'b000000000000;
		12'd1547: color_o = 12'b000000000000;
		12'd1548: color_o = 12'b000000000000;
		12'd1549: color_o = 12'b000000000000;
		12'd1550: color_o = 12'b000000000000;
		12'd1551: color_o = 12'b000000000000;
		12'd1552: color_o = 12'b000000000000;
		12'd1553: color_o = 12'b000000000000;
		12'd1554: color_o = 12'b100000000000;
		12'd1555: color_o = 12'b100000000000;
		12'd1556: color_o = 12'b100000000000;
		12'd1557: color_o = 12'b100000000001;
		12'd1558: color_o = 12'b000000000000;
		12'd1559: color_o = 12'b000011110000;
		12'd1560: color_o = 12'b000011110000;
		12'd1561: color_o = 12'b000011110000;
		12'd1562: color_o = 12'b000011110000;
		12'd1563: color_o = 12'b000011110000;
		12'd1564: color_o = 12'b000011110000;
		12'd1565: color_o = 12'b000011110000;
		12'd1566: color_o = 12'b000011110000;
		12'd1567: color_o = 12'b000011110000;
		12'd1568: color_o = 12'b000011110000;
		12'd1569: color_o = 12'b000011110000;
		12'd1570: color_o = 12'b000000000000;
		12'd1571: color_o = 12'b000000000000;
		12'd1572: color_o = 12'b000000000000;
		12'd1573: color_o = 12'b100000000001;
		12'd1574: color_o = 12'b100000000001;
		12'd1575: color_o = 12'b100000000001;
		12'd1576: color_o = 12'b100000000001;
		12'd1577: color_o = 12'b000000000000;
		12'd1578: color_o = 12'b000000000000;
		12'd1579: color_o = 12'b000000000000;
		12'd1580: color_o = 12'b000000000000;
		12'd1581: color_o = 12'b000000000000;
		12'd1582: color_o = 12'b100000000000;
		12'd1583: color_o = 12'b100000000000;
		12'd1584: color_o = 12'b100000000000;
		12'd1585: color_o = 12'b100000000000;
		12'd1586: color_o = 12'b000000000000;
		12'd1587: color_o = 12'b100000000000;
		12'd1588: color_o = 12'b100000000001;
		12'd1589: color_o = 12'b100000000001;
		12'd1590: color_o = 12'b000000000000;
		12'd1591: color_o = 12'b000011110000;
		12'd1592: color_o = 12'b000011110000;
		12'd1593: color_o = 12'b000011110000;
		12'd1594: color_o = 12'b000011110000;
		12'd1595: color_o = 12'b000011110000;
		12'd1596: color_o = 12'b000011110000;
		12'd1597: color_o = 12'b000011110000;
		12'd1598: color_o = 12'b000011110000;
		12'd1599: color_o = 12'b000011110000;
		12'd1600: color_o = 12'b000011110000;
		12'd1601: color_o = 12'b000000000000;
		12'd1602: color_o = 12'b000000000000;
		12'd1603: color_o = 12'b000000000000;
		12'd1604: color_o = 12'b000000000000;
		12'd1605: color_o = 12'b000000000000;
		12'd1606: color_o = 12'b000000000000;
		12'd1607: color_o = 12'b100000000000;
		12'd1608: color_o = 12'b100000000001;
		12'd1609: color_o = 12'b100000000001;
		12'd1610: color_o = 12'b100000000000;
		12'd1611: color_o = 12'b100000000000;
		12'd1612: color_o = 12'b100000000000;
		12'd1613: color_o = 12'b100000000000;
		12'd1614: color_o = 12'b010000000000;
		12'd1615: color_o = 12'b010000000000;
		12'd1616: color_o = 12'b010000000000;
		12'd1617: color_o = 12'b010000000000;
		12'd1618: color_o = 12'b000000000000;
		12'd1619: color_o = 12'b100000000001;
		12'd1620: color_o = 12'b100000000001;
		12'd1621: color_o = 12'b000000000000;
		12'd1622: color_o = 12'b000000000000;
		12'd1623: color_o = 12'b000011110000;
		12'd1624: color_o = 12'b000011110000;
		12'd1625: color_o = 12'b000011110000;
		12'd1626: color_o = 12'b000011110000;
		12'd1627: color_o = 12'b000011110000;
		12'd1628: color_o = 12'b000011110000;
		12'd1629: color_o = 12'b000011110000;
		12'd1630: color_o = 12'b000011110000;
		12'd1631: color_o = 12'b000011110000;
		12'd1632: color_o = 12'b000011110000;
		12'd1633: color_o = 12'b000000000000;
		12'd1634: color_o = 12'b000000000000;
		12'd1635: color_o = 12'b000000000000;
		12'd1636: color_o = 12'b010000000000;
		12'd1637: color_o = 12'b010000000000;
		12'd1638: color_o = 12'b000000000000;
		12'd1639: color_o = 12'b000000000000;
		12'd1640: color_o = 12'b000000000000;
		12'd1641: color_o = 12'b000000000000;
		12'd1642: color_o = 12'b100000000000;
		12'd1643: color_o = 12'b010000000000;
		12'd1644: color_o = 12'b010000000000;
		12'd1645: color_o = 12'b010000000000;
		12'd1646: color_o = 12'b010000000000;
		12'd1647: color_o = 12'b010000000000;
		12'd1648: color_o = 12'b000000000000;
		12'd1649: color_o = 12'b000000000000;
		12'd1650: color_o = 12'b000000000000;
		12'd1651: color_o = 12'b000000000000;
		12'd1652: color_o = 12'b000000000000;
		12'd1653: color_o = 12'b000000000000;
		12'd1654: color_o = 12'b000000000000;
		12'd1655: color_o = 12'b000011110000;
		12'd1656: color_o = 12'b000011110000;
		12'd1657: color_o = 12'b000011110000;
		12'd1658: color_o = 12'b000011110000;
		12'd1659: color_o = 12'b000011110000;
		12'd1660: color_o = 12'b000011110000;
		12'd1661: color_o = 12'b000011110000;
		12'd1662: color_o = 12'b000011110000;
		12'd1663: color_o = 12'b000011110000;
		12'd1664: color_o = 12'b000011110000;
		12'd1665: color_o = 12'b000000000000;
		12'd1666: color_o = 12'b000000000000;
		12'd1667: color_o = 12'b010000000000;
		12'd1668: color_o = 12'b010000000000;
		12'd1669: color_o = 12'b010000000000;
		12'd1670: color_o = 12'b100000000001;
		12'd1671: color_o = 12'b000000000000;
		12'd1672: color_o = 12'b000000000000;
		12'd1673: color_o = 12'b000000000000;
		12'd1674: color_o = 12'b000000000000;
		12'd1675: color_o = 12'b000000000000;
		12'd1676: color_o = 12'b000000000000;
		12'd1677: color_o = 12'b000000000000;
		12'd1678: color_o = 12'b000000000000;
		12'd1679: color_o = 12'b000000000000;
		12'd1680: color_o = 12'b000000000000;
		12'd1681: color_o = 12'b010000000000;
		12'd1682: color_o = 12'b000000000000;
		12'd1683: color_o = 12'b000000000000;
		12'd1684: color_o = 12'b000000000000;
		12'd1685: color_o = 12'b001000000000;
		12'd1686: color_o = 12'b001000000000;
		12'd1687: color_o = 12'b000000000000;
		12'd1688: color_o = 12'b000011110000;
		12'd1689: color_o = 12'b000011110000;
		12'd1690: color_o = 12'b000011110000;
		12'd1691: color_o = 12'b000011110000;
		12'd1692: color_o = 12'b000011110000;
		12'd1693: color_o = 12'b000011110000;
		12'd1694: color_o = 12'b000011110000;
		12'd1695: color_o = 12'b000011110000;
		12'd1696: color_o = 12'b000011110000;
		12'd1697: color_o = 12'b000000000000;
		12'd1698: color_o = 12'b000000000000;
		12'd1699: color_o = 12'b010000000000;
		12'd1700: color_o = 12'b010000000000;
		12'd1701: color_o = 12'b100000000001;
		12'd1702: color_o = 12'b100000000001;
		12'd1703: color_o = 12'b100000000001;
		12'd1704: color_o = 12'b100000000001;
		12'd1705: color_o = 12'b100000000001;
		12'd1706: color_o = 12'b100000000001;
		12'd1707: color_o = 12'b100000000001;
		12'd1708: color_o = 12'b100000000001;
		12'd1709: color_o = 12'b100000000001;
		12'd1710: color_o = 12'b100000000001;
		12'd1711: color_o = 12'b100000000001;
		12'd1712: color_o = 12'b100000000001;
		12'd1713: color_o = 12'b010000000000;
		12'd1714: color_o = 12'b010000000000;
		12'd1715: color_o = 12'b000000000000;
		12'd1716: color_o = 12'b001000000000;
		12'd1717: color_o = 12'b001000000000;
		12'd1718: color_o = 12'b001000000000;
		12'd1719: color_o = 12'b000000000000;
		12'd1720: color_o = 12'b000011110000;
		12'd1721: color_o = 12'b000011110000;
		12'd1722: color_o = 12'b000011110000;
		12'd1723: color_o = 12'b000011110000;
		12'd1724: color_o = 12'b000011110000;
		12'd1725: color_o = 12'b000011110000;
		12'd1726: color_o = 12'b000011110000;
		12'd1727: color_o = 12'b000011110000;
		12'd1728: color_o = 12'b000011110000;
		12'd1729: color_o = 12'b000000000000;
		12'd1730: color_o = 12'b000000000000;
		12'd1731: color_o = 12'b010000000000;
		12'd1732: color_o = 12'b100000000001;
		12'd1733: color_o = 12'b100000000001;
		12'd1734: color_o = 12'b100000000001;
		12'd1735: color_o = 12'b100000000001;
		12'd1736: color_o = 12'b100000000001;
		12'd1737: color_o = 12'b100000000001;
		12'd1738: color_o = 12'b100000000001;
		12'd1739: color_o = 12'b100000000001;
		12'd1740: color_o = 12'b100000000001;
		12'd1741: color_o = 12'b100000000001;
		12'd1742: color_o = 12'b100000000001;
		12'd1743: color_o = 12'b100000000001;
		12'd1744: color_o = 12'b010000000000;
		12'd1745: color_o = 12'b010000000000;
		12'd1746: color_o = 12'b000000000000;
		12'd1747: color_o = 12'b000000000000;
		12'd1748: color_o = 12'b001000000000;
		12'd1749: color_o = 12'b000000000000;
		12'd1750: color_o = 12'b010000000000;
		12'd1751: color_o = 12'b000000000000;
		12'd1752: color_o = 12'b000011110000;
		12'd1753: color_o = 12'b000011110000;
		12'd1754: color_o = 12'b000011110000;
		12'd1755: color_o = 12'b000011110000;
		12'd1756: color_o = 12'b000011110000;
		12'd1757: color_o = 12'b000011110000;
		12'd1758: color_o = 12'b000011110000;
		12'd1759: color_o = 12'b000011110000;
		12'd1760: color_o = 12'b000011110000;
		12'd1761: color_o = 12'b000000000000;
		12'd1762: color_o = 12'b000000000000;
		12'd1763: color_o = 12'b100000000001;
		12'd1764: color_o = 12'b100000000001;
		12'd1765: color_o = 12'b100000000001;
		12'd1766: color_o = 12'b100000000001;
		12'd1767: color_o = 12'b100000000001;
		12'd1768: color_o = 12'b000000000000;
		12'd1769: color_o = 12'b000000000000;
		12'd1770: color_o = 12'b000000000000;
		12'd1771: color_o = 12'b000000000000;
		12'd1772: color_o = 12'b000000000000;
		12'd1773: color_o = 12'b000000000000;
		12'd1774: color_o = 12'b100000000001;
		12'd1775: color_o = 12'b010000000000;
		12'd1776: color_o = 12'b010000000000;
		12'd1777: color_o = 12'b000000000000;
		12'd1778: color_o = 12'b001000000000;
		12'd1779: color_o = 12'b001000000000;
		12'd1780: color_o = 12'b001000000000;
		12'd1781: color_o = 12'b000000000000;
		12'd1782: color_o = 12'b000000000000;
		12'd1783: color_o = 12'b000000000000;
		12'd1784: color_o = 12'b000011110000;
		12'd1785: color_o = 12'b000011110000;
		12'd1786: color_o = 12'b000011110000;
		12'd1787: color_o = 12'b000011110000;
		12'd1788: color_o = 12'b000011110000;
		12'd1789: color_o = 12'b000011110000;
		12'd1790: color_o = 12'b000011110000;
		12'd1791: color_o = 12'b000011110000;
		12'd1792: color_o = 12'b000011110000;
		12'd1793: color_o = 12'b000000000000;
		12'd1794: color_o = 12'b000000000000;
		12'd1795: color_o = 12'b100000000001;
		12'd1796: color_o = 12'b100000000001;
		12'd1797: color_o = 12'b100000000001;
		12'd1798: color_o = 12'b100000000001;
		12'd1799: color_o = 12'b000000000000;
		12'd1800: color_o = 12'b100000000001;
		12'd1801: color_o = 12'b100000000001;
		12'd1802: color_o = 12'b100000000001;
		12'd1803: color_o = 12'b100000000001;
		12'd1804: color_o = 12'b000000000000;
		12'd1805: color_o = 12'b000000000000;
		12'd1806: color_o = 12'b010000000000;
		12'd1807: color_o = 12'b010000000000;
		12'd1808: color_o = 12'b000000000000;
		12'd1809: color_o = 12'b001000000000;
		12'd1810: color_o = 12'b001000000000;
		12'd1811: color_o = 12'b100000000001;
		12'd1812: color_o = 12'b000000000000;
		12'd1813: color_o = 12'b000000000000;
		12'd1814: color_o = 12'b010000000000;
		12'd1815: color_o = 12'b000000000000;
		12'd1816: color_o = 12'b000011110000;
		12'd1817: color_o = 12'b000011110000;
		12'd1818: color_o = 12'b000011110000;
		12'd1819: color_o = 12'b000011110000;
		12'd1820: color_o = 12'b000011110000;
		12'd1821: color_o = 12'b000011110000;
		12'd1822: color_o = 12'b000011110000;
		12'd1823: color_o = 12'b000011110000;
		12'd1824: color_o = 12'b000011110000;
		12'd1825: color_o = 12'b000011110000;
		12'd1826: color_o = 12'b000000000000;
		12'd1827: color_o = 12'b010000000000;
		12'd1828: color_o = 12'b100000000001;
		12'd1829: color_o = 12'b100000000001;
		12'd1830: color_o = 12'b100000000001;
		12'd1831: color_o = 12'b000000000000;
		12'd1832: color_o = 12'b100000000001;
		12'd1833: color_o = 12'b100000000001;
		12'd1834: color_o = 12'b100000000001;
		12'd1835: color_o = 12'b100000000001;
		12'd1836: color_o = 12'b100000000001;
		12'd1837: color_o = 12'b000000000000;
		12'd1838: color_o = 12'b010000000000;
		12'd1839: color_o = 12'b000000000000;
		12'd1840: color_o = 12'b000000000000;
		12'd1841: color_o = 12'b001000000000;
		12'd1842: color_o = 12'b001000000000;
		12'd1843: color_o = 12'b010000000000;
		12'd1844: color_o = 12'b000000000000;
		12'd1845: color_o = 12'b000000000000;
		12'd1846: color_o = 12'b010000000000;
		12'd1847: color_o = 12'b000000000000;
		12'd1848: color_o = 12'b000000000000;
		12'd1849: color_o = 12'b000011110000;
		12'd1850: color_o = 12'b000011110000;
		12'd1851: color_o = 12'b000011110000;
		12'd1852: color_o = 12'b000011110000;
		12'd1853: color_o = 12'b000011110000;
		12'd1854: color_o = 12'b000011110000;
		12'd1855: color_o = 12'b000011110000;
		12'd1856: color_o = 12'b000011110000;
		12'd1857: color_o = 12'b000011110000;
		12'd1858: color_o = 12'b000000000000;
		12'd1859: color_o = 12'b100000000001;
		12'd1860: color_o = 12'b010000000000;
		12'd1861: color_o = 12'b100000000001;
		12'd1862: color_o = 12'b100000000001;
		12'd1863: color_o = 12'b000000000000;
		12'd1864: color_o = 12'b010000000000;
		12'd1865: color_o = 12'b010000000000;
		12'd1866: color_o = 12'b100000000001;
		12'd1867: color_o = 12'b010000000000;
		12'd1868: color_o = 12'b100000000001;
		12'd1869: color_o = 12'b000000000000;
		12'd1870: color_o = 12'b000000000000;
		12'd1871: color_o = 12'b000000000000;
		12'd1872: color_o = 12'b001000000000;
		12'd1873: color_o = 12'b001000000000;
		12'd1874: color_o = 12'b001000000000;
		12'd1875: color_o = 12'b010000000000;
		12'd1876: color_o = 12'b010000000000;
		12'd1877: color_o = 12'b000000000000;
		12'd1878: color_o = 12'b010000000000;
		12'd1879: color_o = 12'b010000000000;
		12'd1880: color_o = 12'b000000000000;
		12'd1881: color_o = 12'b000011110000;
		12'd1882: color_o = 12'b000011110000;
		12'd1883: color_o = 12'b000011110000;
		12'd1884: color_o = 12'b000011110000;
		12'd1885: color_o = 12'b000011110000;
		12'd1886: color_o = 12'b000011110000;
		12'd1887: color_o = 12'b000011110000;
		12'd1888: color_o = 12'b000011110000;
		12'd1889: color_o = 12'b000000000000;
		12'd1890: color_o = 12'b010000000000;
		12'd1891: color_o = 12'b010000000000;
		12'd1892: color_o = 12'b100000000001;
		12'd1893: color_o = 12'b100000000001;
		12'd1894: color_o = 12'b100000000001;
		12'd1895: color_o = 12'b000000000000;
		12'd1896: color_o = 12'b000000000000;
		12'd1897: color_o = 12'b010000000000;
		12'd1898: color_o = 12'b010000000000;
		12'd1899: color_o = 12'b010000000000;
		12'd1900: color_o = 12'b000000000000;
		12'd1901: color_o = 12'b000000000000;
		12'd1902: color_o = 12'b000000000000;
		12'd1903: color_o = 12'b000000000000;
		12'd1904: color_o = 12'b000000000000;
		12'd1905: color_o = 12'b001000000000;
		12'd1906: color_o = 12'b001000000000;
		12'd1907: color_o = 12'b100000000000;
		12'd1908: color_o = 12'b010000000000;
		12'd1909: color_o = 12'b010000000000;
		12'd1910: color_o = 12'b000000000000;
		12'd1911: color_o = 12'b011000000000;
		12'd1912: color_o = 12'b000000000000;
		12'd1913: color_o = 12'b000011110000;
		12'd1914: color_o = 12'b000011110000;
		12'd1915: color_o = 12'b000011110000;
		12'd1916: color_o = 12'b000011110000;
		12'd1917: color_o = 12'b000011110000;
		12'd1918: color_o = 12'b000011110000;
		12'd1919: color_o = 12'b000011110000;
		12'd1920: color_o = 12'b000011110000;
		12'd1921: color_o = 12'b000000000000;
		12'd1922: color_o = 12'b000000000000;
		12'd1923: color_o = 12'b000000000000;
		12'd1924: color_o = 12'b100000000001;
		12'd1925: color_o = 12'b100000000001;
		12'd1926: color_o = 12'b100000000001;
		12'd1927: color_o = 12'b100000000001;
		12'd1928: color_o = 12'b100000000001;
		12'd1929: color_o = 12'b000000000000;
		12'd1930: color_o = 12'b000000000000;
		12'd1931: color_o = 12'b000000000000;
		12'd1932: color_o = 12'b000000000000;
		12'd1933: color_o = 12'b000011110000;
		12'd1934: color_o = 12'b000000000000;
		12'd1935: color_o = 12'b000000000000;
		12'd1936: color_o = 12'b000000000000;
		12'd1937: color_o = 12'b000000000000;
		12'd1938: color_o = 12'b001000000000;
		12'd1939: color_o = 12'b010000000000;
		12'd1940: color_o = 12'b100000000000;
		12'd1941: color_o = 12'b010000000000;
		12'd1942: color_o = 12'b011000000000;
		12'd1943: color_o = 12'b000000000000;
		12'd1944: color_o = 12'b000000000000;
		12'd1945: color_o = 12'b000011110000;
		12'd1946: color_o = 12'b000011110000;
		12'd1947: color_o = 12'b000011110000;
		12'd1948: color_o = 12'b000011110000;
		12'd1949: color_o = 12'b000011110000;
		12'd1950: color_o = 12'b000011110000;
		12'd1951: color_o = 12'b000011110000;
		12'd1952: color_o = 12'b000011110000;
		12'd1953: color_o = 12'b000000000000;
		12'd1954: color_o = 12'b010000000000;
		12'd1955: color_o = 12'b010000000000;
		12'd1956: color_o = 12'b100000000001;
		12'd1957: color_o = 12'b100000000001;
		12'd1958: color_o = 12'b100000000001;
		12'd1959: color_o = 12'b100000000001;
		12'd1960: color_o = 12'b100000000001;
		12'd1961: color_o = 12'b010000000000;
		12'd1962: color_o = 12'b000000000000;
		12'd1963: color_o = 12'b000011110000;
		12'd1964: color_o = 12'b000011110000;
		12'd1965: color_o = 12'b000011110000;
		12'd1966: color_o = 12'b000011110000;
		12'd1967: color_o = 12'b000000000000;
		12'd1968: color_o = 12'b000000000000;
		12'd1969: color_o = 12'b000000000000;
		12'd1970: color_o = 12'b001000000000;
		12'd1971: color_o = 12'b001000000000;
		12'd1972: color_o = 12'b010000000000;
		12'd1973: color_o = 12'b010000000000;
		12'd1974: color_o = 12'b010000000000;
		12'd1975: color_o = 12'b011000000000;
		12'd1976: color_o = 12'b000000000000;
		12'd1977: color_o = 12'b000000000000;
		12'd1978: color_o = 12'b000011110000;
		12'd1979: color_o = 12'b000011110000;
		12'd1980: color_o = 12'b000011110000;
		12'd1981: color_o = 12'b000011110000;
		12'd1982: color_o = 12'b000011110000;
		12'd1983: color_o = 12'b000011110000;
		12'd1984: color_o = 12'b000011110000;
		12'd1985: color_o = 12'b000000000000;
		12'd1986: color_o = 12'b010000000000;
		12'd1987: color_o = 12'b100000000001;
		12'd1988: color_o = 12'b010000000000;
		12'd1989: color_o = 12'b100000000001;
		12'd1990: color_o = 12'b100000000001;
		12'd1991: color_o = 12'b100000000001;
		12'd1992: color_o = 12'b010000000000;
		12'd1993: color_o = 12'b000000000000;
		12'd1994: color_o = 12'b000011110000;
		12'd1995: color_o = 12'b000011110000;
		12'd1996: color_o = 12'b000011110000;
		12'd1997: color_o = 12'b000011110000;
		12'd1998: color_o = 12'b000011110000;
		12'd1999: color_o = 12'b000011110000;
		12'd2000: color_o = 12'b000000000000;
		12'd2001: color_o = 12'b000000000000;
		12'd2002: color_o = 12'b000000000000;
		12'd2003: color_o = 12'b010000000000;
		12'd2004: color_o = 12'b100000000000;
		12'd2005: color_o = 12'b010000000000;
		12'd2006: color_o = 12'b011000000000;
		12'd2007: color_o = 12'b011000000000;
		12'd2008: color_o = 12'b011000000000;
		12'd2009: color_o = 12'b000000000000;
		12'd2010: color_o = 12'b000000000000;
		12'd2011: color_o = 12'b000011110000;
		12'd2012: color_o = 12'b000011110000;
		12'd2013: color_o = 12'b000011110000;
		12'd2014: color_o = 12'b000011110000;
		12'd2015: color_o = 12'b000011110000;
		12'd2016: color_o = 12'b000011110000;
		12'd2017: color_o = 12'b000000000000;
		12'd2018: color_o = 12'b000000000000;
		12'd2019: color_o = 12'b000000000000;
		12'd2020: color_o = 12'b010000000000;
		12'd2021: color_o = 12'b010000000000;
		12'd2022: color_o = 12'b100000000001;
		12'd2023: color_o = 12'b100000000001;
		12'd2024: color_o = 12'b010000000000;
		12'd2025: color_o = 12'b000000000000;
		12'd2026: color_o = 12'b000000000000;
		12'd2027: color_o = 12'b000000000000;
		12'd2028: color_o = 12'b000011110000;
		12'd2029: color_o = 12'b000011110000;
		12'd2030: color_o = 12'b000011110000;
		12'd2031: color_o = 12'b000011110000;
		12'd2032: color_o = 12'b000011110000;
		12'd2033: color_o = 12'b000000000000;
		12'd2034: color_o = 12'b000000000000;
		12'd2035: color_o = 12'b100000000000;
		12'd2036: color_o = 12'b100000000001;
		12'd2037: color_o = 12'b000000000000;
		12'd2038: color_o = 12'b010000000000;
		12'd2039: color_o = 12'b010000000000;
		12'd2040: color_o = 12'b000000000000;
		12'd2041: color_o = 12'b100000000001;
		12'd2042: color_o = 12'b100000000001;
		12'd2043: color_o = 12'b000000000000;
		12'd2044: color_o = 12'b000000000000;
		12'd2045: color_o = 12'b000000000000;
		12'd2046: color_o = 12'b000011110000;
		12'd2047: color_o = 12'b000011110000;
		12'd2048: color_o = 12'b000000000000;
		12'd2049: color_o = 12'b000000000000;
		12'd2050: color_o = 12'b000000000000;
		12'd2051: color_o = 12'b000000000000;
		12'd2052: color_o = 12'b000000000000;
		12'd2053: color_o = 12'b100000000001;
		12'd2054: color_o = 12'b100000000001;
		12'd2055: color_o = 12'b000000000000;
		12'd2056: color_o = 12'b000000000000;
		12'd2057: color_o = 12'b000000000000;
		12'd2058: color_o = 12'b000000000000;
		12'd2059: color_o = 12'b000000000000;
		12'd2060: color_o = 12'b000011110000;
		12'd2061: color_o = 12'b000011110000;
		12'd2062: color_o = 12'b000011110000;
		12'd2063: color_o = 12'b000011110000;
		12'd2064: color_o = 12'b000011110000;
		12'd2065: color_o = 12'b000000000000;
		12'd2066: color_o = 12'b010000000000;
		12'd2067: color_o = 12'b100000000001;
		12'd2068: color_o = 12'b100000000001;
		12'd2069: color_o = 12'b000000000000;
		12'd2070: color_o = 12'b100000000001;
		12'd2071: color_o = 12'b100000000001;
		12'd2072: color_o = 12'b100000000001;
		12'd2073: color_o = 12'b100000000001;
		12'd2074: color_o = 12'b000000000000;
		12'd2075: color_o = 12'b000000000000;
		12'd2076: color_o = 12'b100000000001;
		12'd2077: color_o = 12'b100000000001;
		12'd2078: color_o = 12'b000000000000;
		12'd2079: color_o = 12'b000011110000;
		12'd2080: color_o = 12'b000000000000;
		12'd2081: color_o = 12'b100000000001;
		12'd2082: color_o = 12'b100000000001;
		12'd2083: color_o = 12'b100000000001;
		12'd2084: color_o = 12'b000000000000;
		12'd2085: color_o = 12'b000000000000;
		12'd2086: color_o = 12'b000000000000;
		12'd2087: color_o = 12'b000000000000;
		12'd2088: color_o = 12'b100000000001;
		12'd2089: color_o = 12'b100000000001;
		12'd2090: color_o = 12'b000000000000;
		12'd2091: color_o = 12'b000000000000;
		12'd2092: color_o = 12'b000000000000;
		12'd2093: color_o = 12'b000011110000;
		12'd2094: color_o = 12'b000011110000;
		12'd2095: color_o = 12'b000011110000;
		12'd2096: color_o = 12'b000011110000;
		12'd2097: color_o = 12'b000000000000;
		12'd2098: color_o = 12'b010000000000;
		12'd2099: color_o = 12'b010000000000;
		12'd2100: color_o = 12'b100000000001;
		12'd2101: color_o = 12'b000000000000;
		12'd2102: color_o = 12'b100000000000;
		12'd2103: color_o = 12'b100000000000;
		12'd2104: color_o = 12'b100000000001;
		12'd2105: color_o = 12'b000000000000;
		12'd2106: color_o = 12'b000000000000;
		12'd2107: color_o = 12'b001000000000;
		12'd2108: color_o = 12'b100000000001;
		12'd2109: color_o = 12'b100000000001;
		12'd2110: color_o = 12'b100000000000;
		12'd2111: color_o = 12'b000000000000;
		12'd2112: color_o = 12'b000000000000;
		12'd2113: color_o = 12'b000000000000;
		12'd2114: color_o = 12'b100000000001;
		12'd2115: color_o = 12'b100000000001;
		12'd2116: color_o = 12'b000000000000;
		12'd2117: color_o = 12'b100000000001;
		12'd2118: color_o = 12'b100000000001;
		12'd2119: color_o = 12'b100000000001;
		12'd2120: color_o = 12'b100000000001;
		12'd2121: color_o = 12'b000000000000;
		12'd2122: color_o = 12'b000000000000;
		12'd2123: color_o = 12'b100000000001;
		12'd2124: color_o = 12'b000000000000;
		12'd2125: color_o = 12'b000000000000;
		12'd2126: color_o = 12'b000011110000;
		12'd2127: color_o = 12'b000011110000;
		12'd2128: color_o = 12'b000000000000;
		12'd2129: color_o = 12'b000000000000;
		12'd2130: color_o = 12'b010000000000;
		12'd2131: color_o = 12'b100000000001;
		12'd2132: color_o = 12'b000000000000;
		12'd2133: color_o = 12'b000000000000;
		12'd2134: color_o = 12'b000000000000;
		12'd2135: color_o = 12'b100000000001;
		12'd2136: color_o = 12'b000000000000;
		12'd2137: color_o = 12'b000000000000;
		12'd2138: color_o = 12'b001000000000;
		12'd2139: color_o = 12'b001000000000;
		12'd2140: color_o = 12'b100000000001;
		12'd2141: color_o = 12'b100000000001;
		12'd2142: color_o = 12'b100000000001;
		12'd2143: color_o = 12'b000000000000;
		12'd2144: color_o = 12'b000011110000;
		12'd2145: color_o = 12'b000000000000;
		12'd2146: color_o = 12'b000000000000;
		12'd2147: color_o = 12'b000000000000;
		12'd2148: color_o = 12'b000000000000;
		12'd2149: color_o = 12'b100000000001;
		12'd2150: color_o = 12'b100000000001;
		12'd2151: color_o = 12'b100000000001;
		12'd2152: color_o = 12'b000000000000;
		12'd2153: color_o = 12'b000000000000;
		12'd2154: color_o = 12'b100000000001;
		12'd2155: color_o = 12'b100000000001;
		12'd2156: color_o = 12'b100000000001;
		12'd2157: color_o = 12'b000000000000;
		12'd2158: color_o = 12'b000000000000;
		12'd2159: color_o = 12'b000000000000;
		12'd2160: color_o = 12'b000000000000;
		12'd2161: color_o = 12'b100000000001;
		12'd2162: color_o = 12'b000000000000;
		12'd2163: color_o = 12'b100000000001;
		12'd2164: color_o = 12'b100000000001;
		12'd2165: color_o = 12'b000000000000;
		12'd2166: color_o = 12'b100000000001;
		12'd2167: color_o = 12'b100000000001;
		12'd2168: color_o = 12'b000000000000;
		12'd2169: color_o = 12'b001000000000;
		12'd2170: color_o = 12'b001000000000;
		12'd2171: color_o = 12'b001000000000;
		12'd2172: color_o = 12'b001000000000;
		12'd2173: color_o = 12'b100000000000;
		12'd2174: color_o = 12'b100000000001;
		12'd2175: color_o = 12'b000000000000;
		12'd2176: color_o = 12'b000011110000;
		12'd2177: color_o = 12'b000011110000;
		12'd2178: color_o = 12'b000000000000;
		12'd2179: color_o = 12'b000000000000;
		12'd2180: color_o = 12'b000000000000;
		12'd2181: color_o = 12'b100000000001;
		12'd2182: color_o = 12'b000000000000;
		12'd2183: color_o = 12'b000000000000;
		12'd2184: color_o = 12'b100000000001;
		12'd2185: color_o = 12'b100000000001;
		12'd2186: color_o = 12'b100000000001;
		12'd2187: color_o = 12'b100000000001;
		12'd2188: color_o = 12'b100000000001;
		12'd2189: color_o = 12'b100000000001;
		12'd2190: color_o = 12'b000000000000;
		12'd2191: color_o = 12'b000000000000;
		12'd2192: color_o = 12'b000000000000;
		12'd2193: color_o = 12'b000000000000;
		12'd2194: color_o = 12'b000000000000;
		12'd2195: color_o = 12'b000000000000;
		12'd2196: color_o = 12'b000000000000;
		12'd2197: color_o = 12'b000000000000;
		12'd2198: color_o = 12'b000000000000;
		12'd2199: color_o = 12'b000000000000;
		12'd2200: color_o = 12'b000000000000;
		12'd2201: color_o = 12'b000000000000;
		12'd2202: color_o = 12'b000000000000;
		12'd2203: color_o = 12'b000000000000;
		12'd2204: color_o = 12'b000000000000;
		12'd2205: color_o = 12'b000000000000;
		12'd2206: color_o = 12'b000000000000;
		12'd2207: color_o = 12'b000000000000;
		12'd2208: color_o = 12'b000011110000;
		12'd2209: color_o = 12'b000011110000;
		12'd2210: color_o = 12'b000011110000;
		12'd2211: color_o = 12'b000000000000;
		12'd2212: color_o = 12'b000000000000;
		12'd2213: color_o = 12'b100000000001;
		12'd2214: color_o = 12'b000000000000;
		12'd2215: color_o = 12'b100000000001;
		12'd2216: color_o = 12'b100000000001;
		12'd2217: color_o = 12'b100000000001;
		12'd2218: color_o = 12'b100000000001;
		12'd2219: color_o = 12'b100000000001;
		12'd2220: color_o = 12'b100000000001;
		12'd2221: color_o = 12'b000000000000;
		12'd2222: color_o = 12'b000000000000;
		12'd2223: color_o = 12'b000011110000;
		12'd2224: color_o = 12'b000011110000;
		12'd2225: color_o = 12'b000011110000;
		12'd2226: color_o = 12'b000011110000;
		12'd2227: color_o = 12'b000011110000;
		12'd2228: color_o = 12'b000011110000;
		12'd2229: color_o = 12'b000000000000;
		12'd2230: color_o = 12'b000000000000;
		12'd2231: color_o = 12'b000000000000;
		12'd2232: color_o = 12'b000000000000;
		12'd2233: color_o = 12'b000011110000;
		12'd2234: color_o = 12'b000011110000;
		12'd2235: color_o = 12'b000011110000;
		12'd2236: color_o = 12'b000011110000;
		12'd2237: color_o = 12'b000011110000;
		12'd2238: color_o = 12'b000011110000;
		12'd2239: color_o = 12'b000011110000;
		12'd2240: color_o = 12'b000011110000;
		12'd2241: color_o = 12'b000011110000;
		12'd2242: color_o = 12'b000011110000;
		12'd2243: color_o = 12'b000011110000;
		12'd2244: color_o = 12'b000000000000;
		12'd2245: color_o = 12'b000000000000;
		12'd2246: color_o = 12'b000000000000;
		12'd2247: color_o = 12'b000000000000;
		12'd2248: color_o = 12'b000000000000;
		12'd2249: color_o = 12'b000000000000;
		12'd2250: color_o = 12'b000000000000;
		12'd2251: color_o = 12'b000000000000;
		12'd2252: color_o = 12'b000000000000;
		12'd2253: color_o = 12'b000000000000;
		12'd2254: color_o = 12'b000011110000;
		12'd2255: color_o = 12'b000011110000;
		12'd2256: color_o = 12'b000011110000;
		12'd2257: color_o = 12'b000011110000;
		12'd2258: color_o = 12'b000011110000;
		12'd2259: color_o = 12'b000011110000;
		12'd2260: color_o = 12'b000011110000;
		12'd2261: color_o = 12'b000011110000;
		12'd2262: color_o = 12'b000011110000;
		12'd2263: color_o = 12'b000011110000;
		12'd2264: color_o = 12'b000011110000;
		12'd2265: color_o = 12'b000011110000;
		12'd2266: color_o = 12'b000011110000;
		12'd2267: color_o = 12'b000011110000;
		12'd2268: color_o = 12'b000011110000;
		12'd2269: color_o = 12'b000011110000;
		12'd2270: color_o = 12'b000011110000;
		12'd2271: color_o = 12'b000011110000;
		12'd2272: color_o = 12'b000011110000;
		12'd2273: color_o = 12'b000011110000;
		12'd2274: color_o = 12'b000011110000;
		12'd2275: color_o = 12'b000011110000;
		12'd2276: color_o = 12'b000011110000;
		12'd2277: color_o = 12'b000011110000;
		12'd2278: color_o = 12'b000011110000;
		12'd2279: color_o = 12'b000011110000;
		12'd2280: color_o = 12'b000011110000;
		12'd2281: color_o = 12'b000011110000;
		12'd2282: color_o = 12'b000011110000;
		12'd2283: color_o = 12'b000011110000;
		12'd2284: color_o = 12'b000011110000;
		12'd2285: color_o = 12'b000011110000;
		12'd2286: color_o = 12'b000011110000;
		12'd2287: color_o = 12'b000011110000;
		12'd2288: color_o = 12'b000011110000;
		12'd2289: color_o = 12'b000011110000;
		12'd2290: color_o = 12'b000011110000;
		12'd2291: color_o = 12'b000011110000;
		12'd2292: color_o = 12'b000011110000;
		12'd2293: color_o = 12'b000011110000;
		12'd2294: color_o = 12'b000011110000;
		12'd2295: color_o = 12'b000011110000;
		12'd2296: color_o = 12'b000011110000;
		12'd2297: color_o = 12'b000011110000;
		12'd2298: color_o = 12'b000011110000;
		12'd2299: color_o = 12'b000011110000;
		12'd2300: color_o = 12'b000011110000;
		12'd2301: color_o = 12'b000011110000;
		12'd2302: color_o = 12'b000011110000;
		12'd2303: color_o = 12'b000011110000;
		12'd2304: color_o = 12'b000011110000;
		12'd2305: color_o = 12'b000000000000;
		12'd2306: color_o = 12'b000000000000;
		12'd2307: color_o = 12'b000000000000;
		12'd2308: color_o = 12'b000000000000;
		12'd2309: color_o = 12'b100000000001;
		12'd2310: color_o = 12'b100000000001;
		12'd2311: color_o = 12'b000000000000;
		12'd2312: color_o = 12'b000000000000;
		12'd2313: color_o = 12'b100000000000;
		12'd2314: color_o = 12'b100000000000;
		12'd2315: color_o = 12'b100000000000;
		12'd2316: color_o = 12'b100000000000;
		12'd2317: color_o = 12'b000000000000;
		12'd2318: color_o = 12'b100000000000;
		12'd2319: color_o = 12'b100000000000;
		12'd2320: color_o = 12'b100000000000;
		12'd2321: color_o = 12'b010000000000;
		12'd2322: color_o = 12'b000000000000;
		12'd2323: color_o = 12'b000000000000;
		12'd2324: color_o = 12'b000011110000;
		12'd2325: color_o = 12'b000011110000;
		12'd2326: color_o = 12'b000011110000;
		12'd2327: color_o = 12'b000011110000;
		12'd2328: color_o = 12'b000011110000;
		12'd2329: color_o = 12'b000011110000;
		12'd2330: color_o = 12'b000011110000;
		12'd2331: color_o = 12'b000011110000;
		12'd2332: color_o = 12'b000011110000;
		12'd2333: color_o = 12'b000011110000;
		12'd2334: color_o = 12'b000011110000;
		12'd2335: color_o = 12'b000011110000;
		12'd2336: color_o = 12'b000011110000;
		12'd2337: color_o = 12'b000000000000;
		12'd2338: color_o = 12'b000000000000;
		12'd2339: color_o = 12'b000000000000;
		12'd2340: color_o = 12'b000000000000;
		12'd2341: color_o = 12'b100000000001;
		12'd2342: color_o = 12'b100000000001;
		12'd2343: color_o = 12'b000000000000;
		12'd2344: color_o = 12'b100000000001;
		12'd2345: color_o = 12'b100000000000;
		12'd2346: color_o = 12'b100000000000;
		12'd2347: color_o = 12'b100000000000;
		12'd2348: color_o = 12'b100000000000;
		12'd2349: color_o = 12'b100000000000;
		12'd2350: color_o = 12'b100000000000;
		12'd2351: color_o = 12'b100000000000;
		12'd2352: color_o = 12'b000000000000;
		12'd2353: color_o = 12'b000000000000;
		12'd2354: color_o = 12'b000000000000;
		12'd2355: color_o = 12'b010000000000;
		12'd2356: color_o = 12'b010000000000;
		12'd2357: color_o = 12'b000000000000;
		12'd2358: color_o = 12'b000011110000;
		12'd2359: color_o = 12'b000011110000;
		12'd2360: color_o = 12'b000011110000;
		12'd2361: color_o = 12'b000011110000;
		12'd2362: color_o = 12'b000011110000;
		12'd2363: color_o = 12'b000011110000;
		12'd2364: color_o = 12'b000011110000;
		12'd2365: color_o = 12'b000011110000;
		12'd2366: color_o = 12'b000011110000;
		12'd2367: color_o = 12'b000011110000;
		12'd2368: color_o = 12'b000011110000;
		12'd2369: color_o = 12'b000000000000;
		12'd2370: color_o = 12'b000000000000;
		12'd2371: color_o = 12'b000000000000;
		12'd2372: color_o = 12'b000000000000;
		12'd2373: color_o = 12'b000000000000;
		12'd2374: color_o = 12'b000000000000;
		12'd2375: color_o = 12'b100000000000;
		12'd2376: color_o = 12'b100000000001;
		12'd2377: color_o = 12'b100000000000;
		12'd2378: color_o = 12'b100000000000;
		12'd2379: color_o = 12'b100000000000;
		12'd2380: color_o = 12'b100000000000;
		12'd2381: color_o = 12'b100000000000;
		12'd2382: color_o = 12'b100000000000;
		12'd2383: color_o = 12'b000000000000;
		12'd2384: color_o = 12'b000000000000;
		12'd2385: color_o = 12'b000000000000;
		12'd2386: color_o = 12'b100000000001;
		12'd2387: color_o = 12'b100000000001;
		12'd2388: color_o = 12'b000000000000;
		12'd2389: color_o = 12'b000000000000;
		12'd2390: color_o = 12'b000011110000;
		12'd2391: color_o = 12'b000011110000;
		12'd2392: color_o = 12'b000011110000;
		12'd2393: color_o = 12'b000011110000;
		12'd2394: color_o = 12'b000011110000;
		12'd2395: color_o = 12'b000011110000;
		12'd2396: color_o = 12'b000011110000;
		12'd2397: color_o = 12'b000011110000;
		12'd2398: color_o = 12'b000011110000;
		12'd2399: color_o = 12'b000011110000;
		12'd2400: color_o = 12'b000011110000;
		12'd2401: color_o = 12'b000011110000;
		12'd2402: color_o = 12'b000000000000;
		12'd2403: color_o = 12'b000000000000;
		12'd2404: color_o = 12'b100000000001;
		12'd2405: color_o = 12'b100000000001;
		12'd2406: color_o = 12'b000000000000;
		12'd2407: color_o = 12'b000000000000;
		12'd2408: color_o = 12'b100000000001;
		12'd2409: color_o = 12'b100000000001;
		12'd2410: color_o = 12'b100000000001;
		12'd2411: color_o = 12'b100000000001;
		12'd2412: color_o = 12'b100000000001;
		12'd2413: color_o = 12'b100000000001;
		12'd2414: color_o = 12'b100000000001;
		12'd2415: color_o = 12'b100000000001;
		12'd2416: color_o = 12'b100000000001;
		12'd2417: color_o = 12'b100000000001;
		12'd2418: color_o = 12'b100000000001;
		12'd2419: color_o = 12'b100000000001;
		12'd2420: color_o = 12'b100000000001;
		12'd2421: color_o = 12'b100000000001;
		12'd2422: color_o = 12'b000000000000;
		12'd2423: color_o = 12'b000011110000;
		12'd2424: color_o = 12'b000011110000;
		12'd2425: color_o = 12'b000011110000;
		12'd2426: color_o = 12'b000011110000;
		12'd2427: color_o = 12'b000011110000;
		12'd2428: color_o = 12'b000011110000;
		12'd2429: color_o = 12'b000011110000;
		12'd2430: color_o = 12'b000011110000;
		12'd2431: color_o = 12'b000011110000;
		12'd2432: color_o = 12'b000011110000;
		12'd2433: color_o = 12'b000011110000;
		12'd2434: color_o = 12'b000000000000;
		12'd2435: color_o = 12'b100000000001;
		12'd2436: color_o = 12'b100000000001;
		12'd2437: color_o = 12'b000000000000;
		12'd2438: color_o = 12'b000000000000;
		12'd2439: color_o = 12'b000000000000;
		12'd2440: color_o = 12'b000000000000;
		12'd2441: color_o = 12'b100000000001;
		12'd2442: color_o = 12'b100000000001;
		12'd2443: color_o = 12'b100000000001;
		12'd2444: color_o = 12'b100000000001;
		12'd2445: color_o = 12'b100000000001;
		12'd2446: color_o = 12'b100000000001;
		12'd2447: color_o = 12'b100000000001;
		12'd2448: color_o = 12'b100000000001;
		12'd2449: color_o = 12'b100000000001;
		12'd2450: color_o = 12'b100000000001;
		12'd2451: color_o = 12'b100000000001;
		12'd2452: color_o = 12'b000000000000;
		12'd2453: color_o = 12'b000000000000;
		12'd2454: color_o = 12'b000000000000;
		12'd2455: color_o = 12'b000000000000;
		12'd2456: color_o = 12'b000011110000;
		12'd2457: color_o = 12'b000011110000;
		12'd2458: color_o = 12'b000011110000;
		12'd2459: color_o = 12'b000011110000;
		12'd2460: color_o = 12'b000011110000;
		12'd2461: color_o = 12'b000011110000;
		12'd2462: color_o = 12'b000011110000;
		12'd2463: color_o = 12'b000011110000;
		12'd2464: color_o = 12'b000011110000;
		12'd2465: color_o = 12'b000011110000;
		12'd2466: color_o = 12'b000000000000;
		12'd2467: color_o = 12'b000000000000;
		12'd2468: color_o = 12'b100000000001;
		12'd2469: color_o = 12'b100000000001;
		12'd2470: color_o = 12'b100000000001;
		12'd2471: color_o = 12'b010000000000;
		12'd2472: color_o = 12'b000000000000;
		12'd2473: color_o = 12'b100000000001;
		12'd2474: color_o = 12'b000000000000;
		12'd2475: color_o = 12'b000000000000;
		12'd2476: color_o = 12'b010000000000;
		12'd2477: color_o = 12'b100000000001;
		12'd2478: color_o = 12'b100000000001;
		12'd2479: color_o = 12'b100000000001;
		12'd2480: color_o = 12'b100000000001;
		12'd2481: color_o = 12'b100000000001;
		12'd2482: color_o = 12'b000000000000;
		12'd2483: color_o = 12'b000000000000;
		12'd2484: color_o = 12'b000000000000;
		12'd2485: color_o = 12'b100000000001;
		12'd2486: color_o = 12'b100000000001;
		12'd2487: color_o = 12'b000000000000;
		12'd2488: color_o = 12'b000011110000;
		12'd2489: color_o = 12'b000011110000;
		12'd2490: color_o = 12'b000011110000;
		12'd2491: color_o = 12'b000011110000;
		12'd2492: color_o = 12'b000011110000;
		12'd2493: color_o = 12'b000011110000;
		12'd2494: color_o = 12'b000011110000;
		12'd2495: color_o = 12'b000011110000;
		12'd2496: color_o = 12'b000011110000;
		12'd2497: color_o = 12'b000011110000;
		12'd2498: color_o = 12'b000000000000;
		12'd2499: color_o = 12'b000000000000;
		12'd2500: color_o = 12'b100000000001;
		12'd2501: color_o = 12'b100000000001;
		12'd2502: color_o = 12'b100000000001;
		12'd2503: color_o = 12'b000000000000;
		12'd2504: color_o = 12'b000000000000;
		12'd2505: color_o = 12'b100000000001;
		12'd2506: color_o = 12'b010000000000;
		12'd2507: color_o = 12'b000000000000;
		12'd2508: color_o = 12'b010000000000;
		12'd2509: color_o = 12'b100000000001;
		12'd2510: color_o = 12'b010000000000;
		12'd2511: color_o = 12'b100000000001;
		12'd2512: color_o = 12'b100000000001;
		12'd2513: color_o = 12'b100000000001;
		12'd2514: color_o = 12'b100000000001;
		12'd2515: color_o = 12'b100000000001;
		12'd2516: color_o = 12'b100000000001;
		12'd2517: color_o = 12'b100000000001;
		12'd2518: color_o = 12'b100000000001;
		12'd2519: color_o = 12'b100000000001;
		12'd2520: color_o = 12'b000000000000;
		12'd2521: color_o = 12'b000011110000;
		12'd2522: color_o = 12'b000011110000;
		12'd2523: color_o = 12'b000011110000;
		12'd2524: color_o = 12'b000011110000;
		12'd2525: color_o = 12'b000011110000;
		12'd2526: color_o = 12'b000011110000;
		12'd2527: color_o = 12'b000011110000;
		12'd2528: color_o = 12'b000011110000;
		12'd2529: color_o = 12'b000011110000;
		12'd2530: color_o = 12'b000000000000;
		12'd2531: color_o = 12'b000000000000;
		12'd2532: color_o = 12'b000000000000;
		12'd2533: color_o = 12'b100000000001;
		12'd2534: color_o = 12'b100000000001;
		12'd2535: color_o = 12'b000000000000;
		12'd2536: color_o = 12'b000000000000;
		12'd2537: color_o = 12'b100000000001;
		12'd2538: color_o = 12'b010000000000;
		12'd2539: color_o = 12'b000000000000;
		12'd2540: color_o = 12'b100000000001;
		12'd2541: color_o = 12'b010000000000;
		12'd2542: color_o = 12'b100000000001;
		12'd2543: color_o = 12'b010000000000;
		12'd2544: color_o = 12'b100000000001;
		12'd2545: color_o = 12'b100000000001;
		12'd2546: color_o = 12'b000000000000;
		12'd2547: color_o = 12'b100000000001;
		12'd2548: color_o = 12'b100000000001;
		12'd2549: color_o = 12'b100000000001;
		12'd2550: color_o = 12'b100000000001;
		12'd2551: color_o = 12'b100000000001;
		12'd2552: color_o = 12'b000000000000;
		12'd2553: color_o = 12'b000011110000;
		12'd2554: color_o = 12'b000011110000;
		12'd2555: color_o = 12'b000011110000;
		12'd2556: color_o = 12'b000011110000;
		12'd2557: color_o = 12'b000011110000;
		12'd2558: color_o = 12'b000011110000;
		12'd2559: color_o = 12'b000011110000;
		12'd2560: color_o = 12'b000011110000;
		12'd2561: color_o = 12'b000011110000;
		12'd2562: color_o = 12'b000011110000;
		12'd2563: color_o = 12'b000000000000;
		12'd2564: color_o = 12'b000000000000;
		12'd2565: color_o = 12'b000000000000;
		12'd2566: color_o = 12'b000000000000;
		12'd2567: color_o = 12'b000000000000;
		12'd2568: color_o = 12'b000000000000;
		12'd2569: color_o = 12'b000000000000;
		12'd2570: color_o = 12'b000000000000;
		12'd2571: color_o = 12'b000000000000;
		12'd2572: color_o = 12'b000000000000;
		12'd2573: color_o = 12'b100000000001;
		12'd2574: color_o = 12'b010000000000;
		12'd2575: color_o = 12'b100000000001;
		12'd2576: color_o = 12'b010000000000;
		12'd2577: color_o = 12'b100000000001;
		12'd2578: color_o = 12'b000000000000;
		12'd2579: color_o = 12'b100000000001;
		12'd2580: color_o = 12'b100000000001;
		12'd2581: color_o = 12'b100000000001;
		12'd2582: color_o = 12'b100000000001;
		12'd2583: color_o = 12'b100000000001;
		12'd2584: color_o = 12'b000000000000;
		12'd2585: color_o = 12'b000011110000;
		12'd2586: color_o = 12'b000011110000;
		12'd2587: color_o = 12'b000011110000;
		12'd2588: color_o = 12'b000011110000;
		12'd2589: color_o = 12'b000011110000;
		12'd2590: color_o = 12'b000011110000;
		12'd2591: color_o = 12'b000011110000;
		12'd2592: color_o = 12'b000011110000;
		12'd2593: color_o = 12'b000011110000;
		12'd2594: color_o = 12'b000011110000;
		12'd2595: color_o = 12'b000000000000;
		12'd2596: color_o = 12'b000000000000;
		12'd2597: color_o = 12'b000000000000;
		12'd2598: color_o = 12'b000000000000;
		12'd2599: color_o = 12'b000000000000;
		12'd2600: color_o = 12'b000000000000;
		12'd2601: color_o = 12'b000000000000;
		12'd2602: color_o = 12'b000000000000;
		12'd2603: color_o = 12'b000000000000;
		12'd2604: color_o = 12'b000000000000;
		12'd2605: color_o = 12'b000000000000;
		12'd2606: color_o = 12'b000000000000;
		12'd2607: color_o = 12'b010000000000;
		12'd2608: color_o = 12'b010000000000;
		12'd2609: color_o = 12'b100000000001;
		12'd2610: color_o = 12'b000000000000;
		12'd2611: color_o = 12'b010000000000;
		12'd2612: color_o = 12'b100000000001;
		12'd2613: color_o = 12'b100000000001;
		12'd2614: color_o = 12'b010000000000;
		12'd2615: color_o = 12'b000000000000;
		12'd2616: color_o = 12'b000000000000;
		12'd2617: color_o = 12'b000011110000;
		12'd2618: color_o = 12'b000011110000;
		12'd2619: color_o = 12'b000011110000;
		12'd2620: color_o = 12'b000011110000;
		12'd2621: color_o = 12'b000011110000;
		12'd2622: color_o = 12'b000011110000;
		12'd2623: color_o = 12'b000011110000;
		12'd2624: color_o = 12'b000011110000;
		12'd2625: color_o = 12'b000011110000;
		12'd2626: color_o = 12'b000011110000;
		12'd2627: color_o = 12'b000000000000;
		12'd2628: color_o = 12'b000000000000;
		12'd2629: color_o = 12'b000000000000;
		12'd2630: color_o = 12'b000000000000;
		12'd2631: color_o = 12'b010000000000;
		12'd2632: color_o = 12'b010000000000;
		12'd2633: color_o = 12'b010000000000;
		12'd2634: color_o = 12'b000000000000;
		12'd2635: color_o = 12'b000000000000;
		12'd2636: color_o = 12'b000000000000;
		12'd2637: color_o = 12'b000000000000;
		12'd2638: color_o = 12'b000000000000;
		12'd2639: color_o = 12'b000000000000;
		12'd2640: color_o = 12'b000000000000;
		12'd2641: color_o = 12'b100000000001;
		12'd2642: color_o = 12'b000000000000;
		12'd2643: color_o = 12'b000000000000;
		12'd2644: color_o = 12'b010000000000;
		12'd2645: color_o = 12'b010000000000;
		12'd2646: color_o = 12'b010000000000;
		12'd2647: color_o = 12'b000000000000;
		12'd2648: color_o = 12'b000011110000;
		12'd2649: color_o = 12'b000011110000;
		12'd2650: color_o = 12'b000011110000;
		12'd2651: color_o = 12'b000011110000;
		12'd2652: color_o = 12'b000011110000;
		12'd2653: color_o = 12'b000011110000;
		12'd2654: color_o = 12'b000011110000;
		12'd2655: color_o = 12'b000011110000;
		12'd2656: color_o = 12'b000011110000;
		12'd2657: color_o = 12'b000011110000;
		12'd2658: color_o = 12'b000000000000;
		12'd2659: color_o = 12'b000000000000;
		12'd2660: color_o = 12'b000000000000;
		12'd2661: color_o = 12'b000000000000;
		12'd2662: color_o = 12'b010000000000;
		12'd2663: color_o = 12'b010000000000;
		12'd2664: color_o = 12'b010000000000;
		12'd2665: color_o = 12'b010000000000;
		12'd2666: color_o = 12'b010000000000;
		12'd2667: color_o = 12'b000000000000;
		12'd2668: color_o = 12'b000000000000;
		12'd2669: color_o = 12'b000011110000;
		12'd2670: color_o = 12'b000000000000;
		12'd2671: color_o = 12'b000000000000;
		12'd2672: color_o = 12'b100000000001;
		12'd2673: color_o = 12'b100000000001;
		12'd2674: color_o = 12'b100000000001;
		12'd2675: color_o = 12'b100000000001;
		12'd2676: color_o = 12'b000000000000;
		12'd2677: color_o = 12'b000000000000;
		12'd2678: color_o = 12'b000000000000;
		12'd2679: color_o = 12'b000000000000;
		12'd2680: color_o = 12'b000011110000;
		12'd2681: color_o = 12'b000011110000;
		12'd2682: color_o = 12'b000011110000;
		12'd2683: color_o = 12'b000011110000;
		12'd2684: color_o = 12'b000011110000;
		12'd2685: color_o = 12'b000011110000;
		12'd2686: color_o = 12'b000011110000;
		12'd2687: color_o = 12'b000011110000;
		12'd2688: color_o = 12'b000011110000;
		12'd2689: color_o = 12'b000011110000;
		12'd2690: color_o = 12'b000000000000;
		12'd2691: color_o = 12'b000000000000;
		12'd2692: color_o = 12'b000000000000;
		12'd2693: color_o = 12'b010000000000;
		12'd2694: color_o = 12'b010000000000;
		12'd2695: color_o = 12'b000000000000;
		12'd2696: color_o = 12'b010000000000;
		12'd2697: color_o = 12'b010000000000;
		12'd2698: color_o = 12'b000000000000;
		12'd2699: color_o = 12'b000000000000;
		12'd2700: color_o = 12'b000011110000;
		12'd2701: color_o = 12'b000011110000;
		12'd2702: color_o = 12'b000000000000;
		12'd2703: color_o = 12'b000000000000;
		12'd2704: color_o = 12'b100000000001;
		12'd2705: color_o = 12'b100000000001;
		12'd2706: color_o = 12'b100000000001;
		12'd2707: color_o = 12'b100000000001;
		12'd2708: color_o = 12'b100000000001;
		12'd2709: color_o = 12'b100000000001;
		12'd2710: color_o = 12'b000000000000;
		12'd2711: color_o = 12'b000000000000;
		12'd2712: color_o = 12'b000000000000;
		12'd2713: color_o = 12'b000011110000;
		12'd2714: color_o = 12'b000011110000;
		12'd2715: color_o = 12'b000011110000;
		12'd2716: color_o = 12'b000011110000;
		12'd2717: color_o = 12'b000011110000;
		12'd2718: color_o = 12'b000011110000;
		12'd2719: color_o = 12'b000011110000;
		12'd2720: color_o = 12'b000011110000;
		12'd2721: color_o = 12'b000011110000;
		12'd2722: color_o = 12'b000000000000;
		12'd2723: color_o = 12'b000000000000;
		12'd2724: color_o = 12'b000000000000;
		12'd2725: color_o = 12'b000000000000;
		12'd2726: color_o = 12'b000000000000;
		12'd2727: color_o = 12'b000000000000;
		12'd2728: color_o = 12'b000000000000;
		12'd2729: color_o = 12'b000000000000;
		12'd2730: color_o = 12'b000000000000;
		12'd2731: color_o = 12'b000000000000;
		12'd2732: color_o = 12'b000011110000;
		12'd2733: color_o = 12'b000011110000;
		12'd2734: color_o = 12'b000011110000;
		12'd2735: color_o = 12'b000000000000;
		12'd2736: color_o = 12'b000000000000;
		12'd2737: color_o = 12'b000000000000;
		12'd2738: color_o = 12'b100000000001;
		12'd2739: color_o = 12'b100000000001;
		12'd2740: color_o = 12'b100000000001;
		12'd2741: color_o = 12'b000000000000;
		12'd2742: color_o = 12'b000000000000;
		12'd2743: color_o = 12'b000000000000;
		12'd2744: color_o = 12'b000000000000;
		12'd2745: color_o = 12'b000000000000;
		12'd2746: color_o = 12'b000011110000;
		12'd2747: color_o = 12'b000011110000;
		12'd2748: color_o = 12'b000011110000;
		12'd2749: color_o = 12'b000011110000;
		12'd2750: color_o = 12'b000011110000;
		12'd2751: color_o = 12'b000011110000;
		12'd2752: color_o = 12'b000011110000;
		12'd2753: color_o = 12'b000011110000;
		12'd2754: color_o = 12'b000000000000;
		12'd2755: color_o = 12'b000000000000;
		12'd2756: color_o = 12'b000000000000;
		12'd2757: color_o = 12'b010000000000;
		12'd2758: color_o = 12'b000000000000;
		12'd2759: color_o = 12'b000000000000;
		12'd2760: color_o = 12'b000000000000;
		12'd2761: color_o = 12'b010000000000;
		12'd2762: color_o = 12'b000000000000;
		12'd2763: color_o = 12'b000011110000;
		12'd2764: color_o = 12'b000011110000;
		12'd2765: color_o = 12'b000011110000;
		12'd2766: color_o = 12'b000011110000;
		12'd2767: color_o = 12'b000000000000;
		12'd2768: color_o = 12'b000000000000;
		12'd2769: color_o = 12'b000000000000;
		12'd2770: color_o = 12'b000000000000;
		12'd2771: color_o = 12'b000000000000;
		12'd2772: color_o = 12'b000000000000;
		12'd2773: color_o = 12'b000000000000;
		12'd2774: color_o = 12'b000000000000;
		12'd2775: color_o = 12'b100000000001;
		12'd2776: color_o = 12'b100000000001;
		12'd2777: color_o = 12'b000000000000;
		12'd2778: color_o = 12'b000000000000;
		12'd2779: color_o = 12'b000011110000;
		12'd2780: color_o = 12'b000011110000;
		12'd2781: color_o = 12'b000011110000;
		12'd2782: color_o = 12'b000011110000;
		12'd2783: color_o = 12'b000011110000;
		12'd2784: color_o = 12'b000011110000;
		12'd2785: color_o = 12'b000000000000;
		12'd2786: color_o = 12'b000000000000;
		12'd2787: color_o = 12'b000000000000;
		12'd2788: color_o = 12'b010000000000;
		12'd2789: color_o = 12'b000000000000;
		12'd2790: color_o = 12'b010000000000;
		12'd2791: color_o = 12'b000000000000;
		12'd2792: color_o = 12'b000000000000;
		12'd2793: color_o = 12'b010000000000;
		12'd2794: color_o = 12'b000011110000;
		12'd2795: color_o = 12'b000011110000;
		12'd2796: color_o = 12'b000011110000;
		12'd2797: color_o = 12'b000011110000;
		12'd2798: color_o = 12'b000011110000;
		12'd2799: color_o = 12'b000000000000;
		12'd2800: color_o = 12'b100000000001;
		12'd2801: color_o = 12'b100000000001;
		12'd2802: color_o = 12'b100000000001;
		12'd2803: color_o = 12'b000000000000;
		12'd2804: color_o = 12'b100000000001;
		12'd2805: color_o = 12'b100000000001;
		12'd2806: color_o = 12'b100000000001;
		12'd2807: color_o = 12'b100000000001;
		12'd2808: color_o = 12'b000000000000;
		12'd2809: color_o = 12'b000000000000;
		12'd2810: color_o = 12'b000000000000;
		12'd2811: color_o = 12'b000000000000;
		12'd2812: color_o = 12'b000011110000;
		12'd2813: color_o = 12'b000011110000;
		12'd2814: color_o = 12'b000011110000;
		12'd2815: color_o = 12'b000011110000;
		12'd2816: color_o = 12'b000011110000;
		12'd2817: color_o = 12'b000000000000;
		12'd2818: color_o = 12'b000000000000;
		12'd2819: color_o = 12'b000000000000;
		12'd2820: color_o = 12'b000000000000;
		12'd2821: color_o = 12'b010000000000;
		12'd2822: color_o = 12'b000000000000;
		12'd2823: color_o = 12'b000000000000;
		12'd2824: color_o = 12'b000000000000;
		12'd2825: color_o = 12'b010000000000;
		12'd2826: color_o = 12'b000000000000;
		12'd2827: color_o = 12'b000011110000;
		12'd2828: color_o = 12'b000011110000;
		12'd2829: color_o = 12'b000011110000;
		12'd2830: color_o = 12'b000011110000;
		12'd2831: color_o = 12'b000000000000;
		12'd2832: color_o = 12'b100000000001;
		12'd2833: color_o = 12'b100000000001;
		12'd2834: color_o = 12'b100000000001;
		12'd2835: color_o = 12'b000000000000;
		12'd2836: color_o = 12'b100000000001;
		12'd2837: color_o = 12'b100000000001;
		12'd2838: color_o = 12'b100000000001;
		12'd2839: color_o = 12'b000000000000;
		12'd2840: color_o = 12'b000000000000;
		12'd2841: color_o = 12'b100000000001;
		12'd2842: color_o = 12'b100000000001;
		12'd2843: color_o = 12'b000000000000;
		12'd2844: color_o = 12'b000000000000;
		12'd2845: color_o = 12'b000011110000;
		12'd2846: color_o = 12'b000011110000;
		12'd2847: color_o = 12'b000011110000;
		12'd2848: color_o = 12'b000000000000;
		12'd2849: color_o = 12'b000000000000;
		12'd2850: color_o = 12'b000000000000;
		12'd2851: color_o = 12'b000000000000;
		12'd2852: color_o = 12'b010000000000;
		12'd2853: color_o = 12'b000000000000;
		12'd2854: color_o = 12'b100000000001;
		12'd2855: color_o = 12'b100000000001;
		12'd2856: color_o = 12'b100000000001;
		12'd2857: color_o = 12'b100000000001;
		12'd2858: color_o = 12'b000000000000;
		12'd2859: color_o = 12'b000011110000;
		12'd2860: color_o = 12'b000011110000;
		12'd2861: color_o = 12'b000000000000;
		12'd2862: color_o = 12'b000000000000;
		12'd2863: color_o = 12'b000000000000;
		12'd2864: color_o = 12'b010000000000;
		12'd2865: color_o = 12'b100000000001;
		12'd2866: color_o = 12'b000000000000;
		12'd2867: color_o = 12'b000000000000;
		12'd2868: color_o = 12'b000000000000;
		12'd2869: color_o = 12'b100000000001;
		12'd2870: color_o = 12'b000000000000;
		12'd2871: color_o = 12'b000000000000;
		12'd2872: color_o = 12'b100000000001;
		12'd2873: color_o = 12'b100000000001;
		12'd2874: color_o = 12'b100000000001;
		12'd2875: color_o = 12'b100000000001;
		12'd2876: color_o = 12'b000000000000;
		12'd2877: color_o = 12'b000000000000;
		12'd2878: color_o = 12'b000011110000;
		12'd2879: color_o = 12'b000011110000;
		12'd2880: color_o = 12'b000011110000;
		12'd2881: color_o = 12'b000000000000;
		12'd2882: color_o = 12'b000000000000;
		12'd2883: color_o = 12'b000000000000;
		12'd2884: color_o = 12'b000000000000;
		12'd2885: color_o = 12'b000000000000;
		12'd2886: color_o = 12'b000000000000;
		12'd2887: color_o = 12'b000000000000;
		12'd2888: color_o = 12'b000000000000;
		12'd2889: color_o = 12'b000000000000;
		12'd2890: color_o = 12'b000000000000;
		12'd2891: color_o = 12'b000011110000;
		12'd2892: color_o = 12'b000011110000;
		12'd2893: color_o = 12'b000011110000;
		12'd2894: color_o = 12'b000000000000;
		12'd2895: color_o = 12'b000000000000;
		12'd2896: color_o = 12'b000000000000;
		12'd2897: color_o = 12'b100000000001;
		12'd2898: color_o = 12'b100000000001;
		12'd2899: color_o = 12'b000000000000;
		12'd2900: color_o = 12'b000000000000;
		12'd2901: color_o = 12'b100000000001;
		12'd2902: color_o = 12'b000000000000;
		12'd2903: color_o = 12'b010000000000;
		12'd2904: color_o = 12'b010000000000;
		12'd2905: color_o = 12'b100000000001;
		12'd2906: color_o = 12'b100000000001;
		12'd2907: color_o = 12'b100000000001;
		12'd2908: color_o = 12'b100000000001;
		12'd2909: color_o = 12'b000000000000;
		12'd2910: color_o = 12'b000011110000;
		12'd2911: color_o = 12'b000011110000;
		12'd2912: color_o = 12'b000011110000;
		12'd2913: color_o = 12'b000011110000;
		12'd2914: color_o = 12'b000000000000;
		12'd2915: color_o = 12'b000000000000;
		12'd2916: color_o = 12'b000000000000;
		12'd2917: color_o = 12'b000000000000;
		12'd2918: color_o = 12'b000000000000;
		12'd2919: color_o = 12'b010000000000;
		12'd2920: color_o = 12'b100000000001;
		12'd2921: color_o = 12'b010000000000;
		12'd2922: color_o = 12'b000000000000;
		12'd2923: color_o = 12'b000000000000;
		12'd2924: color_o = 12'b000011110000;
		12'd2925: color_o = 12'b000011110000;
		12'd2926: color_o = 12'b000011110000;
		12'd2927: color_o = 12'b000011110000;
		12'd2928: color_o = 12'b000000000000;
		12'd2929: color_o = 12'b000000000000;
		12'd2930: color_o = 12'b000000000000;
		12'd2931: color_o = 12'b000000000000;
		12'd2932: color_o = 12'b000000000000;
		12'd2933: color_o = 12'b000000000000;
		12'd2934: color_o = 12'b000000000000;
		12'd2935: color_o = 12'b000000000000;
		12'd2936: color_o = 12'b010000000000;
		12'd2937: color_o = 12'b100000000001;
		12'd2938: color_o = 12'b100000000001;
		12'd2939: color_o = 12'b100000000001;
		12'd2940: color_o = 12'b100000000001;
		12'd2941: color_o = 12'b000000000000;
		12'd2942: color_o = 12'b000011110000;
		12'd2943: color_o = 12'b000011110000;
		12'd2944: color_o = 12'b000011110000;
		12'd2945: color_o = 12'b000011110000;
		12'd2946: color_o = 12'b000011110000;
		12'd2947: color_o = 12'b000000000000;
		12'd2948: color_o = 12'b000000000000;
		12'd2949: color_o = 12'b000000000000;
		12'd2950: color_o = 12'b000000000000;
		12'd2951: color_o = 12'b000000000000;
		12'd2952: color_o = 12'b100000000001;
		12'd2953: color_o = 12'b010000000000;
		12'd2954: color_o = 12'b010000000000;
		12'd2955: color_o = 12'b000000000000;
		12'd2956: color_o = 12'b000000000000;
		12'd2957: color_o = 12'b000011110000;
		12'd2958: color_o = 12'b000011110000;
		12'd2959: color_o = 12'b000011110000;
		12'd2960: color_o = 12'b000011110000;
		12'd2961: color_o = 12'b000011110000;
		12'd2962: color_o = 12'b000011110000;
		12'd2963: color_o = 12'b000000000000;
		12'd2964: color_o = 12'b000000000000;
		12'd2965: color_o = 12'b000000000000;
		12'd2966: color_o = 12'b000000000000;
		12'd2967: color_o = 12'b000000000000;
		12'd2968: color_o = 12'b000000000000;
		12'd2969: color_o = 12'b100000000001;
		12'd2970: color_o = 12'b100000000001;
		12'd2971: color_o = 12'b100000000001;
		12'd2972: color_o = 12'b100000000001;
		12'd2973: color_o = 12'b000000000000;
		12'd2974: color_o = 12'b000011110000;
		12'd2975: color_o = 12'b000011110000;
		12'd2976: color_o = 12'b000011110000;
		12'd2977: color_o = 12'b000011110000;
		12'd2978: color_o = 12'b000011110000;
		12'd2979: color_o = 12'b000011110000;
		12'd2980: color_o = 12'b000011110000;
		12'd2981: color_o = 12'b000000000000;
		12'd2982: color_o = 12'b000000000000;
		12'd2983: color_o = 12'b000000000000;
		12'd2984: color_o = 12'b000000000000;
		12'd2985: color_o = 12'b000000000000;
		12'd2986: color_o = 12'b000000000000;
		12'd2987: color_o = 12'b000000000000;
		12'd2988: color_o = 12'b000000000000;
		12'd2989: color_o = 12'b000000000000;
		12'd2990: color_o = 12'b000011110000;
		12'd2991: color_o = 12'b000011110000;
		12'd2992: color_o = 12'b000011110000;
		12'd2993: color_o = 12'b000011110000;
		12'd2994: color_o = 12'b000011110000;
		12'd2995: color_o = 12'b000011110000;
		12'd2996: color_o = 12'b000011110000;
		12'd2997: color_o = 12'b000011110000;
		12'd2998: color_o = 12'b000011110000;
		12'd2999: color_o = 12'b000000000000;
		12'd3000: color_o = 12'b000000000000;
		12'd3001: color_o = 12'b000000000000;
		12'd3002: color_o = 12'b000000000000;
		12'd3003: color_o = 12'b000000000000;
		12'd3004: color_o = 12'b000000000000;
		12'd3005: color_o = 12'b000000000000;
		12'd3006: color_o = 12'b000011110000;
		12'd3007: color_o = 12'b000011110000;
		12'd3008: color_o = 12'b000011110000;
		12'd3009: color_o = 12'b000011110000;
		12'd3010: color_o = 12'b000011110000;
		12'd3011: color_o = 12'b000011110000;
		12'd3012: color_o = 12'b000011110000;
		12'd3013: color_o = 12'b000011110000;
		12'd3014: color_o = 12'b000000000000;
		12'd3015: color_o = 12'b000000000000;
		12'd3016: color_o = 12'b000000000000;
		12'd3017: color_o = 12'b000000000000;
		12'd3018: color_o = 12'b000000000000;
		12'd3019: color_o = 12'b000000000000;
		12'd3020: color_o = 12'b000000000000;
		12'd3021: color_o = 12'b000000000000;
		12'd3022: color_o = 12'b000011110000;
		12'd3023: color_o = 12'b000011110000;
		12'd3024: color_o = 12'b000011110000;
		12'd3025: color_o = 12'b000011110000;
		12'd3026: color_o = 12'b000011110000;
		12'd3027: color_o = 12'b000011110000;
		12'd3028: color_o = 12'b000011110000;
		12'd3029: color_o = 12'b000011110000;
		12'd3030: color_o = 12'b000011110000;
		12'd3031: color_o = 12'b000011110000;
		12'd3032: color_o = 12'b000011110000;
		12'd3033: color_o = 12'b000011110000;
		12'd3034: color_o = 12'b000011110000;
		12'd3035: color_o = 12'b000011110000;
		12'd3036: color_o = 12'b000011110000;
		12'd3037: color_o = 12'b000011110000;
		12'd3038: color_o = 12'b000011110000;
		12'd3039: color_o = 12'b000011110000;
		12'd3040: color_o = 12'b000011110000;
		12'd3041: color_o = 12'b000011110000;
		12'd3042: color_o = 12'b000011110000;
		12'd3043: color_o = 12'b000011110000;
		12'd3044: color_o = 12'b000011110000;
		12'd3045: color_o = 12'b000011110000;
		12'd3046: color_o = 12'b000011110000;
		12'd3047: color_o = 12'b000000000000;
		12'd3048: color_o = 12'b000000000000;
		12'd3049: color_o = 12'b000000000000;
		12'd3050: color_o = 12'b000000000000;
		12'd3051: color_o = 12'b000000000000;
		12'd3052: color_o = 12'b000000000000;
		12'd3053: color_o = 12'b000000000000;
		12'd3054: color_o = 12'b000011110000;
		12'd3055: color_o = 12'b000011110000;
		12'd3056: color_o = 12'b000011110000;
		12'd3057: color_o = 12'b000011110000;
		12'd3058: color_o = 12'b000011110000;
		12'd3059: color_o = 12'b000011110000;
		12'd3060: color_o = 12'b000011110000;
		12'd3061: color_o = 12'b000011110000;
		12'd3062: color_o = 12'b000011110000;
		12'd3063: color_o = 12'b000011110000;
		12'd3064: color_o = 12'b000011110000;
		12'd3065: color_o = 12'b000011110000;
		12'd3066: color_o = 12'b000011110000;
		12'd3067: color_o = 12'b000011110000;
		12'd3068: color_o = 12'b000011110000;
		12'd3069: color_o = 12'b000011110000;
		12'd3070: color_o = 12'b000011110000;
		12'd3071: color_o = 12'b000011110000;

        default: color_o = 12'h000;
    endcase       
    
endmodule
