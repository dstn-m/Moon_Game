`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/12/2023 09:28:42 PM
// Design Name: 
// Module Name: char_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module char_rom(
    input clk_i,
    input [12:0] addr,
    output reg [11:0] color_o
    );

reg[12:0] addr_in;

always @ (posedge clk_i) begin
    addr_in <= addr;            // latch in current address
end    
    
always @*
    case(addr_in)
		13'd0: color_o = 12'b000011110000;
		13'd1: color_o = 12'b000011110000;
		13'd2: color_o = 12'b000011110000;
		13'd3: color_o = 12'b000011110000;
		13'd4: color_o = 12'b000011110000;
		13'd5: color_o = 12'b000011110000;
		13'd6: color_o = 12'b000011110000;
		13'd7: color_o = 12'b000011110000;
		13'd8: color_o = 12'b000011110000;
		13'd9: color_o = 12'b000011110000;
		13'd10: color_o = 12'b000011110000;
		13'd11: color_o = 12'b000011110000;
		13'd12: color_o = 12'b000011110000;
		13'd13: color_o = 12'b000011110000;
		13'd14: color_o = 12'b000011110000;
		13'd15: color_o = 12'b000011110000;
		13'd16: color_o = 12'b000011110000;
		13'd17: color_o = 12'b000011110000;
		13'd18: color_o = 12'b000011110000;
		13'd19: color_o = 12'b000011110000;
		13'd20: color_o = 12'b000011110000;
		13'd21: color_o = 12'b000011110000;
		13'd22: color_o = 12'b000011110000;
		13'd23: color_o = 12'b000011110000;
		13'd24: color_o = 12'b000011110000;
		13'd25: color_o = 12'b000011110000;
		13'd26: color_o = 12'b000011110000;
		13'd27: color_o = 12'b000011110000;
		13'd28: color_o = 12'b000011110000;
		13'd29: color_o = 12'b000011110000;
		13'd30: color_o = 12'b000011110000;
		13'd31: color_o = 12'b000011110000;
		13'd32: color_o = 12'b000011110000;
		13'd33: color_o = 12'b000011110000;
		13'd34: color_o = 12'b000011110000;
		13'd35: color_o = 12'b000011110000;
		13'd36: color_o = 12'b000011110000;
		13'd37: color_o = 12'b000011110000;
		13'd38: color_o = 12'b000011110000;
		13'd39: color_o = 12'b000011110000;
		13'd40: color_o = 12'b000011110000;
		13'd41: color_o = 12'b000011110000;
		13'd42: color_o = 12'b000011110000;
		13'd43: color_o = 12'b000011110000;
		13'd44: color_o = 12'b000011110000;
		13'd45: color_o = 12'b000011110000;
		13'd46: color_o = 12'b000011110000;
		13'd47: color_o = 12'b000011110000;
		13'd48: color_o = 12'b000011110000;
		13'd49: color_o = 12'b000011110000;
		13'd50: color_o = 12'b000011110000;
		13'd51: color_o = 12'b000011110000;
		13'd52: color_o = 12'b000011110000;
		13'd53: color_o = 12'b000011110000;
		13'd54: color_o = 12'b000011110000;
		13'd55: color_o = 12'b000011110000;
		13'd56: color_o = 12'b000011110000;
		13'd57: color_o = 12'b000011110000;
		13'd58: color_o = 12'b000011110000;
		13'd59: color_o = 12'b000011110000;
		13'd60: color_o = 12'b000011110000;
		13'd61: color_o = 12'b000011110000;
		13'd62: color_o = 12'b000011110000;
		13'd63: color_o = 12'b000011110000;
		13'd64: color_o = 12'b000011110000;
		13'd65: color_o = 12'b000011110000;
		13'd66: color_o = 12'b000011110000;
		13'd67: color_o = 12'b000011110000;
		13'd68: color_o = 12'b000011110000;
		13'd69: color_o = 12'b000011110000;
		13'd70: color_o = 12'b000011110000;
		13'd71: color_o = 12'b000011110000;
		13'd72: color_o = 12'b000011110000;
		13'd73: color_o = 12'b000011110000;
		13'd74: color_o = 12'b000011110000;
		13'd75: color_o = 12'b000011110000;
		13'd76: color_o = 12'b000011110000;
		13'd77: color_o = 12'b000011110000;
		13'd78: color_o = 12'b000000000000;
		13'd79: color_o = 12'b000000000000;
		13'd80: color_o = 12'b000000000000;
		13'd81: color_o = 12'b011000000000;
		13'd82: color_o = 12'b011000000000;
		13'd83: color_o = 12'b011000000000;
		13'd84: color_o = 12'b000011110000;
		13'd85: color_o = 12'b000011110000;
		13'd86: color_o = 12'b000011110000;
		13'd87: color_o = 12'b000011110000;
		13'd88: color_o = 12'b000011110000;
		13'd89: color_o = 12'b000011110000;
		13'd90: color_o = 12'b000011110000;
		13'd91: color_o = 12'b000011110000;
		13'd92: color_o = 12'b000011110000;
		13'd93: color_o = 12'b000011110000;
		13'd94: color_o = 12'b000011110000;
		13'd95: color_o = 12'b000011110000;
		13'd96: color_o = 12'b000011110000;
		13'd97: color_o = 12'b000011110000;
		13'd98: color_o = 12'b000011110000;
		13'd99: color_o = 12'b000011110000;
		13'd100: color_o = 12'b000011110000;
		13'd101: color_o = 12'b000011110000;
		13'd102: color_o = 12'b000011110000;
		13'd103: color_o = 12'b000011110000;
		13'd104: color_o = 12'b000011110000;
		13'd105: color_o = 12'b000011110000;
		13'd106: color_o = 12'b000011110000;
		13'd107: color_o = 12'b000011110000;
		13'd108: color_o = 12'b000011110000;
		13'd109: color_o = 12'b000011110000;
		13'd110: color_o = 12'b000011110000;
		13'd111: color_o = 12'b000011110000;
		13'd112: color_o = 12'b000011110000;
		13'd113: color_o = 12'b000011110000;
		13'd114: color_o = 12'b000011110000;
		13'd115: color_o = 12'b000011110000;
		13'd116: color_o = 12'b000011110000;
		13'd117: color_o = 12'b000011110000;
		13'd118: color_o = 12'b000011110000;
		13'd119: color_o = 12'b000011110000;
		13'd120: color_o = 12'b000011110000;
		13'd121: color_o = 12'b000011110000;
		13'd122: color_o = 12'b000011110000;
		13'd123: color_o = 12'b000011110000;
		13'd124: color_o = 12'b000011110000;
		13'd125: color_o = 12'b000011110000;
		13'd126: color_o = 12'b000011110000;
		13'd127: color_o = 12'b000011110000;
		13'd128: color_o = 12'b000011110000;
		13'd129: color_o = 12'b000011110000;
		13'd130: color_o = 12'b000011110000;
		13'd131: color_o = 12'b000011110000;
		13'd132: color_o = 12'b000011110000;
		13'd133: color_o = 12'b000011110000;
		13'd134: color_o = 12'b000011110000;
		13'd135: color_o = 12'b000011110000;
		13'd136: color_o = 12'b000011110000;
		13'd137: color_o = 12'b000011110000;
		13'd138: color_o = 12'b000011110000;
		13'd139: color_o = 12'b000011110000;
		13'd140: color_o = 12'b000011110000;
		13'd141: color_o = 12'b000000000000;
		13'd142: color_o = 12'b000000000000;
		13'd143: color_o = 12'b000000000000;
		13'd144: color_o = 12'b100000000000;
		13'd145: color_o = 12'b011000000000;
		13'd146: color_o = 12'b011000000000;
		13'd147: color_o = 12'b011000000000;
		13'd148: color_o = 12'b011000000000;
		13'd149: color_o = 12'b011000000000;
		13'd150: color_o = 12'b011000000000;
		13'd151: color_o = 12'b011000000000;
		13'd152: color_o = 12'b000011110000;
		13'd153: color_o = 12'b000011110000;
		13'd154: color_o = 12'b000011110000;
		13'd155: color_o = 12'b000011110000;
		13'd156: color_o = 12'b000011110000;
		13'd157: color_o = 12'b000011110000;
		13'd158: color_o = 12'b000011110000;
		13'd159: color_o = 12'b000011110000;
		13'd160: color_o = 12'b000011110000;
		13'd161: color_o = 12'b000011110000;
		13'd162: color_o = 12'b000011110000;
		13'd163: color_o = 12'b000011110000;
		13'd164: color_o = 12'b000011110000;
		13'd165: color_o = 12'b000011110000;
		13'd166: color_o = 12'b000011110000;
		13'd167: color_o = 12'b000011110000;
		13'd168: color_o = 12'b000011110000;
		13'd169: color_o = 12'b000011110000;
		13'd170: color_o = 12'b000011110000;
		13'd171: color_o = 12'b000011110000;
		13'd172: color_o = 12'b000011110000;
		13'd173: color_o = 12'b000011110000;
		13'd174: color_o = 12'b000011110000;
		13'd175: color_o = 12'b000011110000;
		13'd176: color_o = 12'b000011110000;
		13'd177: color_o = 12'b000011110000;
		13'd178: color_o = 12'b000011110000;
		13'd179: color_o = 12'b000011110000;
		13'd180: color_o = 12'b000011110000;
		13'd181: color_o = 12'b000011110000;
		13'd182: color_o = 12'b000011110000;
		13'd183: color_o = 12'b000011110000;
		13'd184: color_o = 12'b000011110000;
		13'd185: color_o = 12'b000011110000;
		13'd186: color_o = 12'b000011110000;
		13'd187: color_o = 12'b000011110000;
		13'd188: color_o = 12'b000011110000;
		13'd189: color_o = 12'b000011110000;
		13'd190: color_o = 12'b000011110000;
		13'd191: color_o = 12'b000011110000;
		13'd192: color_o = 12'b000011110000;
		13'd193: color_o = 12'b000011110000;
		13'd194: color_o = 12'b000011110000;
		13'd195: color_o = 12'b000011110000;
		13'd196: color_o = 12'b000011110000;
		13'd197: color_o = 12'b000011110000;
		13'd198: color_o = 12'b000011110000;
		13'd199: color_o = 12'b000011110000;
		13'd200: color_o = 12'b000011110000;
		13'd201: color_o = 12'b000011110000;
		13'd202: color_o = 12'b000011110000;
		13'd203: color_o = 12'b000000000000;
		13'd204: color_o = 12'b000000000000;
		13'd205: color_o = 12'b000000000000;
		13'd206: color_o = 12'b100000000000;
		13'd207: color_o = 12'b100000000000;
		13'd208: color_o = 12'b100000000000;
		13'd209: color_o = 12'b100000000000;
		13'd210: color_o = 12'b100000000000;
		13'd211: color_o = 12'b100000000000;
		13'd212: color_o = 12'b011000000000;
		13'd213: color_o = 12'b011000000000;
		13'd214: color_o = 12'b100000000000;
		13'd215: color_o = 12'b011000000000;
		13'd216: color_o = 12'b011000000000;
		13'd217: color_o = 12'b011000000000;
		13'd218: color_o = 12'b011000000000;
		13'd219: color_o = 12'b011000000000;
		13'd220: color_o = 12'b011000000000;
		13'd221: color_o = 12'b000011110000;
		13'd222: color_o = 12'b000011110000;
		13'd223: color_o = 12'b000011110000;
		13'd224: color_o = 12'b000011110000;
		13'd225: color_o = 12'b000011110000;
		13'd226: color_o = 12'b000011110000;
		13'd227: color_o = 12'b000011110000;
		13'd228: color_o = 12'b000011110000;
		13'd229: color_o = 12'b000011110000;
		13'd230: color_o = 12'b000011110000;
		13'd231: color_o = 12'b000011110000;
		13'd232: color_o = 12'b000011110000;
		13'd233: color_o = 12'b000011110000;
		13'd234: color_o = 12'b000011110000;
		13'd235: color_o = 12'b000011110000;
		13'd236: color_o = 12'b000011110000;
		13'd237: color_o = 12'b000011110000;
		13'd238: color_o = 12'b000011110000;
		13'd239: color_o = 12'b000011110000;
		13'd240: color_o = 12'b000011110000;
		13'd241: color_o = 12'b000011110000;
		13'd242: color_o = 12'b000011110000;
		13'd243: color_o = 12'b000011110000;
		13'd244: color_o = 12'b000011110000;
		13'd245: color_o = 12'b000011110000;
		13'd246: color_o = 12'b000011110000;
		13'd247: color_o = 12'b000011110000;
		13'd248: color_o = 12'b000011110000;
		13'd249: color_o = 12'b000011110000;
		13'd250: color_o = 12'b000011110000;
		13'd251: color_o = 12'b000011110000;
		13'd252: color_o = 12'b000011110000;
		13'd253: color_o = 12'b000011110000;
		13'd254: color_o = 12'b000011110000;
		13'd255: color_o = 12'b000011110000;
		13'd256: color_o = 12'b000011110000;
		13'd257: color_o = 12'b000011110000;
		13'd258: color_o = 12'b000011110000;
		13'd259: color_o = 12'b000011110000;
		13'd260: color_o = 12'b000011110000;
		13'd261: color_o = 12'b000011110000;
		13'd262: color_o = 12'b000011110000;
		13'd263: color_o = 12'b000011110000;
		13'd264: color_o = 12'b000011110000;
		13'd265: color_o = 12'b000011110000;
		13'd266: color_o = 12'b000000000000;
		13'd267: color_o = 12'b000000000000;
		13'd268: color_o = 12'b000000000000;
		13'd269: color_o = 12'b000000000000;
		13'd270: color_o = 12'b100000000000;
		13'd271: color_o = 12'b100000000000;
		13'd272: color_o = 12'b100000000000;
		13'd273: color_o = 12'b100000000000;
		13'd274: color_o = 12'b100000000000;
		13'd275: color_o = 12'b100000000000;
		13'd276: color_o = 12'b100000000000;
		13'd277: color_o = 12'b100000000000;
		13'd278: color_o = 12'b100000000000;
		13'd279: color_o = 12'b100000000000;
		13'd280: color_o = 12'b100000000000;
		13'd281: color_o = 12'b100000000000;
		13'd282: color_o = 12'b011000000000;
		13'd283: color_o = 12'b011000000000;
		13'd284: color_o = 12'b011000000000;
		13'd285: color_o = 12'b011000000000;
		13'd286: color_o = 12'b011000000000;
		13'd287: color_o = 12'b000011110000;
		13'd288: color_o = 12'b000011110000;
		13'd289: color_o = 12'b000011110000;
		13'd290: color_o = 12'b000011110000;
		13'd291: color_o = 12'b000011110000;
		13'd292: color_o = 12'b000011110000;
		13'd293: color_o = 12'b000011110000;
		13'd294: color_o = 12'b000011110000;
		13'd295: color_o = 12'b000011110000;
		13'd296: color_o = 12'b000011110000;
		13'd297: color_o = 12'b000011110000;
		13'd298: color_o = 12'b000011110000;
		13'd299: color_o = 12'b000011110000;
		13'd300: color_o = 12'b000011110000;
		13'd301: color_o = 12'b000011110000;
		13'd302: color_o = 12'b000011110000;
		13'd303: color_o = 12'b000011110000;
		13'd304: color_o = 12'b000011110000;
		13'd305: color_o = 12'b000011110000;
		13'd306: color_o = 12'b000011110000;
		13'd307: color_o = 12'b000011110000;
		13'd308: color_o = 12'b000011110000;
		13'd309: color_o = 12'b000011110000;
		13'd310: color_o = 12'b000011110000;
		13'd311: color_o = 12'b000011110000;
		13'd312: color_o = 12'b000011110000;
		13'd313: color_o = 12'b000011110000;
		13'd314: color_o = 12'b000011110000;
		13'd315: color_o = 12'b000011110000;
		13'd316: color_o = 12'b000011110000;
		13'd317: color_o = 12'b000011110000;
		13'd318: color_o = 12'b000011110000;
		13'd319: color_o = 12'b000011110000;
		13'd320: color_o = 12'b000011110000;
		13'd321: color_o = 12'b000011110000;
		13'd322: color_o = 12'b000011110000;
		13'd323: color_o = 12'b000011110000;
		13'd324: color_o = 12'b000011110000;
		13'd325: color_o = 12'b000011110000;
		13'd326: color_o = 12'b000011110000;
		13'd327: color_o = 12'b000011110000;
		13'd328: color_o = 12'b000011110000;
		13'd329: color_o = 12'b000000000000;
		13'd330: color_o = 12'b000000000000;
		13'd331: color_o = 12'b100001000000;
		13'd332: color_o = 12'b000000000000;
		13'd333: color_o = 12'b000000000000;
		13'd334: color_o = 12'b000000000000;
		13'd335: color_o = 12'b000000000000;
		13'd336: color_o = 12'b100000000000;
		13'd337: color_o = 12'b100000000000;
		13'd338: color_o = 12'b100000000000;
		13'd339: color_o = 12'b100000000000;
		13'd340: color_o = 12'b100000000000;
		13'd341: color_o = 12'b100000000000;
		13'd342: color_o = 12'b011000000000;
		13'd343: color_o = 12'b011000000000;
		13'd344: color_o = 12'b011000000000;
		13'd345: color_o = 12'b100000000000;
		13'd346: color_o = 12'b100000000000;
		13'd347: color_o = 12'b100000000000;
		13'd348: color_o = 12'b011000000000;
		13'd349: color_o = 12'b011000000000;
		13'd350: color_o = 12'b011000000000;
		13'd351: color_o = 12'b011000000000;
		13'd352: color_o = 12'b000011110000;
		13'd353: color_o = 12'b000011110000;
		13'd354: color_o = 12'b000011110000;
		13'd355: color_o = 12'b000011110000;
		13'd356: color_o = 12'b000011110000;
		13'd357: color_o = 12'b000011110000;
		13'd358: color_o = 12'b000011110000;
		13'd359: color_o = 12'b000011110000;
		13'd360: color_o = 12'b000011110000;
		13'd361: color_o = 12'b000011110000;
		13'd362: color_o = 12'b000011110000;
		13'd363: color_o = 12'b000011110000;
		13'd364: color_o = 12'b000011110000;
		13'd365: color_o = 12'b000011110000;
		13'd366: color_o = 12'b000011110000;
		13'd367: color_o = 12'b000011110000;
		13'd368: color_o = 12'b000011110000;
		13'd369: color_o = 12'b000011110000;
		13'd370: color_o = 12'b000011110000;
		13'd371: color_o = 12'b000011110000;
		13'd372: color_o = 12'b000011110000;
		13'd373: color_o = 12'b000011110000;
		13'd374: color_o = 12'b000011110000;
		13'd375: color_o = 12'b000011110000;
		13'd376: color_o = 12'b000011110000;
		13'd377: color_o = 12'b000011110000;
		13'd378: color_o = 12'b000011110000;
		13'd379: color_o = 12'b000011110000;
		13'd380: color_o = 12'b000011110000;
		13'd381: color_o = 12'b000011110000;
		13'd382: color_o = 12'b000011110000;
		13'd383: color_o = 12'b000011110000;
		13'd384: color_o = 12'b000011110000;
		13'd385: color_o = 12'b000011110000;
		13'd386: color_o = 12'b000011110000;
		13'd387: color_o = 12'b000011110000;
		13'd388: color_o = 12'b000011110000;
		13'd389: color_o = 12'b000011110000;
		13'd390: color_o = 12'b000011110000;
		13'd391: color_o = 12'b000011110000;
		13'd392: color_o = 12'b100001000000;
		13'd393: color_o = 12'b100001000000;
		13'd394: color_o = 12'b100001000000;
		13'd395: color_o = 12'b000000000000;
		13'd396: color_o = 12'b000000000000;
		13'd397: color_o = 12'b100000000001;
		13'd398: color_o = 12'b100000000001;
		13'd399: color_o = 12'b100000000001;
		13'd400: color_o = 12'b100000000001;
		13'd401: color_o = 12'b000000000000;
		13'd402: color_o = 12'b000000000000;
		13'd403: color_o = 12'b000000000000;
		13'd404: color_o = 12'b100000000000;
		13'd405: color_o = 12'b100000000000;
		13'd406: color_o = 12'b100000000000;
		13'd407: color_o = 12'b100000000000;
		13'd408: color_o = 12'b100000000000;
		13'd409: color_o = 12'b100000000000;
		13'd410: color_o = 12'b011000000000;
		13'd411: color_o = 12'b011000000000;
		13'd412: color_o = 12'b011000000000;
		13'd413: color_o = 12'b011000000000;
		13'd414: color_o = 12'b100000000000;
		13'd415: color_o = 12'b100000000000;
		13'd416: color_o = 12'b100000000000;
		13'd417: color_o = 12'b000011110000;
		13'd418: color_o = 12'b000011110000;
		13'd419: color_o = 12'b000011110000;
		13'd420: color_o = 12'b000011110000;
		13'd421: color_o = 12'b000011110000;
		13'd422: color_o = 12'b000011110000;
		13'd423: color_o = 12'b000011110000;
		13'd424: color_o = 12'b000011110000;
		13'd425: color_o = 12'b000011110000;
		13'd426: color_o = 12'b000011110000;
		13'd427: color_o = 12'b000011110000;
		13'd428: color_o = 12'b000011110000;
		13'd429: color_o = 12'b000011110000;
		13'd430: color_o = 12'b000011110000;
		13'd431: color_o = 12'b000011110000;
		13'd432: color_o = 12'b000011110000;
		13'd433: color_o = 12'b000011110000;
		13'd434: color_o = 12'b000011110000;
		13'd435: color_o = 12'b000011110000;
		13'd436: color_o = 12'b000011110000;
		13'd437: color_o = 12'b000011110000;
		13'd438: color_o = 12'b000011110000;
		13'd439: color_o = 12'b000011110000;
		13'd440: color_o = 12'b000011110000;
		13'd441: color_o = 12'b000011110000;
		13'd442: color_o = 12'b000011110000;
		13'd443: color_o = 12'b000011110000;
		13'd444: color_o = 12'b000011110000;
		13'd445: color_o = 12'b000011110000;
		13'd446: color_o = 12'b000011110000;
		13'd447: color_o = 12'b000011110000;
		13'd448: color_o = 12'b000011110000;
		13'd449: color_o = 12'b000011110000;
		13'd450: color_o = 12'b000011110000;
		13'd451: color_o = 12'b000011110000;
		13'd452: color_o = 12'b000011110000;
		13'd453: color_o = 12'b000011110000;
		13'd454: color_o = 12'b000011110000;
		13'd455: color_o = 12'b000011110000;
		13'd456: color_o = 12'b100001000000;
		13'd457: color_o = 12'b100001000000;
		13'd458: color_o = 12'b000000000000;
		13'd459: color_o = 12'b000000000000;
		13'd460: color_o = 12'b100000000001;
		13'd461: color_o = 12'b100000000001;
		13'd462: color_o = 12'b100000000001;
		13'd463: color_o = 12'b100000000001;
		13'd464: color_o = 12'b100000000001;
		13'd465: color_o = 12'b100000000001;
		13'd466: color_o = 12'b100000000001;
		13'd467: color_o = 12'b000000000000;
		13'd468: color_o = 12'b000000000000;
		13'd469: color_o = 12'b000000000000;
		13'd470: color_o = 12'b000000000000;
		13'd471: color_o = 12'b000000000000;
		13'd472: color_o = 12'b000000000000;
		13'd473: color_o = 12'b100000000000;
		13'd474: color_o = 12'b100000000000;
		13'd475: color_o = 12'b100000000000;
		13'd476: color_o = 12'b100000000000;
		13'd477: color_o = 12'b100000000000;
		13'd478: color_o = 12'b100000000000;
		13'd479: color_o = 12'b100000000000;
		13'd480: color_o = 12'b100000000000;
		13'd481: color_o = 12'b000011110000;
		13'd482: color_o = 12'b000011110000;
		13'd483: color_o = 12'b000011110000;
		13'd484: color_o = 12'b000011110000;
		13'd485: color_o = 12'b000011110000;
		13'd486: color_o = 12'b000011110000;
		13'd487: color_o = 12'b000011110000;
		13'd488: color_o = 12'b000011110000;
		13'd489: color_o = 12'b000011110000;
		13'd490: color_o = 12'b000011110000;
		13'd491: color_o = 12'b000011110000;
		13'd492: color_o = 12'b000011110000;
		13'd493: color_o = 12'b000011110000;
		13'd494: color_o = 12'b000011110000;
		13'd495: color_o = 12'b000011110000;
		13'd496: color_o = 12'b000011110000;
		13'd497: color_o = 12'b000011110000;
		13'd498: color_o = 12'b000011110000;
		13'd499: color_o = 12'b000011110000;
		13'd500: color_o = 12'b000011110000;
		13'd501: color_o = 12'b000011110000;
		13'd502: color_o = 12'b000011110000;
		13'd503: color_o = 12'b000011110000;
		13'd504: color_o = 12'b000011110000;
		13'd505: color_o = 12'b000011110000;
		13'd506: color_o = 12'b000011110000;
		13'd507: color_o = 12'b000011110000;
		13'd508: color_o = 12'b000011110000;
		13'd509: color_o = 12'b000011110000;
		13'd510: color_o = 12'b000011110000;
		13'd511: color_o = 12'b000011110000;
		13'd512: color_o = 12'b000011110000;
		13'd513: color_o = 12'b000011110000;
		13'd514: color_o = 12'b000011110000;
		13'd515: color_o = 12'b000011110000;
		13'd516: color_o = 12'b000011110000;
		13'd517: color_o = 12'b000011110000;
		13'd518: color_o = 12'b000011110000;
		13'd519: color_o = 12'b000011110000;
		13'd520: color_o = 12'b000000000000;
		13'd521: color_o = 12'b000000000000;
		13'd522: color_o = 12'b000000000000;
		13'd523: color_o = 12'b100000000001;
		13'd524: color_o = 12'b100000000001;
		13'd525: color_o = 12'b100000000001;
		13'd526: color_o = 12'b100000000001;
		13'd527: color_o = 12'b100000000001;
		13'd528: color_o = 12'b100000000001;
		13'd529: color_o = 12'b000000000000;
		13'd530: color_o = 12'b000000000000;
		13'd531: color_o = 12'b000000000000;
		13'd532: color_o = 12'b000000000000;
		13'd533: color_o = 12'b000000000000;
		13'd534: color_o = 12'b100000000001;
		13'd535: color_o = 12'b100000000001;
		13'd536: color_o = 12'b000000000000;
		13'd537: color_o = 12'b000000000000;
		13'd538: color_o = 12'b100000000000;
		13'd539: color_o = 12'b100000000000;
		13'd540: color_o = 12'b100000000000;
		13'd541: color_o = 12'b100000000000;
		13'd542: color_o = 12'b100000000000;
		13'd543: color_o = 12'b100000000000;
		13'd544: color_o = 12'b100000000000;
		13'd545: color_o = 12'b000011110000;
		13'd546: color_o = 12'b000011110000;
		13'd547: color_o = 12'b000011110000;
		13'd548: color_o = 12'b000011110000;
		13'd549: color_o = 12'b000011110000;
		13'd550: color_o = 12'b000011110000;
		13'd551: color_o = 12'b000011110000;
		13'd552: color_o = 12'b000011110000;
		13'd553: color_o = 12'b000011110000;
		13'd554: color_o = 12'b000011110000;
		13'd555: color_o = 12'b000011110000;
		13'd556: color_o = 12'b000011110000;
		13'd557: color_o = 12'b000011110000;
		13'd558: color_o = 12'b000011110000;
		13'd559: color_o = 12'b000011110000;
		13'd560: color_o = 12'b000011110000;
		13'd561: color_o = 12'b000011110000;
		13'd562: color_o = 12'b000011110000;
		13'd563: color_o = 12'b000011110000;
		13'd564: color_o = 12'b000011110000;
		13'd565: color_o = 12'b000011110000;
		13'd566: color_o = 12'b000011110000;
		13'd567: color_o = 12'b000011110000;
		13'd568: color_o = 12'b000011110000;
		13'd569: color_o = 12'b000011110000;
		13'd570: color_o = 12'b000011110000;
		13'd571: color_o = 12'b000011110000;
		13'd572: color_o = 12'b000011110000;
		13'd573: color_o = 12'b000011110000;
		13'd574: color_o = 12'b000011110000;
		13'd575: color_o = 12'b000011110000;
		13'd576: color_o = 12'b000011110000;
		13'd577: color_o = 12'b000011110000;
		13'd578: color_o = 12'b000011110000;
		13'd579: color_o = 12'b000011110000;
		13'd580: color_o = 12'b000011110000;
		13'd581: color_o = 12'b000011110000;
		13'd582: color_o = 12'b000011110000;
		13'd583: color_o = 12'b000011110000;
		13'd584: color_o = 12'b000000000000;
		13'd585: color_o = 12'b000000000000;
		13'd586: color_o = 12'b100000000001;
		13'd587: color_o = 12'b100000000001;
		13'd588: color_o = 12'b100000000001;
		13'd589: color_o = 12'b000000000000;
		13'd590: color_o = 12'b000000000000;
		13'd591: color_o = 12'b000000000000;
		13'd592: color_o = 12'b000000000000;
		13'd593: color_o = 12'b000000000000;
		13'd594: color_o = 12'b100000000001;
		13'd595: color_o = 12'b100000000001;
		13'd596: color_o = 12'b100000000001;
		13'd597: color_o = 12'b100000000001;
		13'd598: color_o = 12'b100000000001;
		13'd599: color_o = 12'b100000000001;
		13'd600: color_o = 12'b100000000001;
		13'd601: color_o = 12'b000000000000;
		13'd602: color_o = 12'b000000000000;
		13'd603: color_o = 12'b000000000000;
		13'd604: color_o = 12'b000000000000;
		13'd605: color_o = 12'b000000000000;
		13'd606: color_o = 12'b000000000000;
		13'd607: color_o = 12'b000000000000;
		13'd608: color_o = 12'b000000000000;
		13'd609: color_o = 12'b111000010010;
		13'd610: color_o = 12'b000011110000;
		13'd611: color_o = 12'b000011110000;
		13'd612: color_o = 12'b000011110000;
		13'd613: color_o = 12'b000011110000;
		13'd614: color_o = 12'b000011110000;
		13'd615: color_o = 12'b000011110000;
		13'd616: color_o = 12'b000011110000;
		13'd617: color_o = 12'b000011110000;
		13'd618: color_o = 12'b000011110000;
		13'd619: color_o = 12'b000011110000;
		13'd620: color_o = 12'b000011110000;
		13'd621: color_o = 12'b000011110000;
		13'd622: color_o = 12'b000011110000;
		13'd623: color_o = 12'b000011110000;
		13'd624: color_o = 12'b000011110000;
		13'd625: color_o = 12'b000011110000;
		13'd626: color_o = 12'b000011110000;
		13'd627: color_o = 12'b000011110000;
		13'd628: color_o = 12'b000011110000;
		13'd629: color_o = 12'b000011110000;
		13'd630: color_o = 12'b000011110000;
		13'd631: color_o = 12'b000011110000;
		13'd632: color_o = 12'b000011110000;
		13'd633: color_o = 12'b000011110000;
		13'd634: color_o = 12'b000011110000;
		13'd635: color_o = 12'b000011110000;
		13'd636: color_o = 12'b000011110000;
		13'd637: color_o = 12'b000011110000;
		13'd638: color_o = 12'b000011110000;
		13'd639: color_o = 12'b000011110000;
		13'd640: color_o = 12'b000011110000;
		13'd641: color_o = 12'b000011110000;
		13'd642: color_o = 12'b000011110000;
		13'd643: color_o = 12'b000011110000;
		13'd644: color_o = 12'b000011110000;
		13'd645: color_o = 12'b000011110000;
		13'd646: color_o = 12'b000011110000;
		13'd647: color_o = 12'b000011110000;
		13'd648: color_o = 12'b000000000000;
		13'd649: color_o = 12'b000000000000;
		13'd650: color_o = 12'b100000000001;
		13'd651: color_o = 12'b000000000000;
		13'd652: color_o = 12'b000000000000;
		13'd653: color_o = 12'b000000000000;
		13'd654: color_o = 12'b100001000000;
		13'd655: color_o = 12'b100001000000;
		13'd656: color_o = 12'b000000000000;
		13'd657: color_o = 12'b100000000001;
		13'd658: color_o = 12'b100000000001;
		13'd659: color_o = 12'b100000000001;
		13'd660: color_o = 12'b000000000000;
		13'd661: color_o = 12'b000000000000;
		13'd662: color_o = 12'b000000000000;
		13'd663: color_o = 12'b000000000000;
		13'd664: color_o = 12'b000000000000;
		13'd665: color_o = 12'b111000010010;
		13'd666: color_o = 12'b111000010010;
		13'd667: color_o = 12'b111000010010;
		13'd668: color_o = 12'b111000010010;
		13'd669: color_o = 12'b111000010010;
		13'd670: color_o = 12'b111000010010;
		13'd671: color_o = 12'b111000010010;
		13'd672: color_o = 12'b111000010010;
		13'd673: color_o = 12'b111000010010;
		13'd674: color_o = 12'b111000010010;
		13'd675: color_o = 12'b000011110000;
		13'd676: color_o = 12'b000011110000;
		13'd677: color_o = 12'b000011110000;
		13'd678: color_o = 12'b000011110000;
		13'd679: color_o = 12'b000011110000;
		13'd680: color_o = 12'b000011110000;
		13'd681: color_o = 12'b000011110000;
		13'd682: color_o = 12'b000011110000;
		13'd683: color_o = 12'b000011110000;
		13'd684: color_o = 12'b000011110000;
		13'd685: color_o = 12'b000011110000;
		13'd686: color_o = 12'b000011110000;
		13'd687: color_o = 12'b000011110000;
		13'd688: color_o = 12'b000011110000;
		13'd689: color_o = 12'b000011110000;
		13'd690: color_o = 12'b000011110000;
		13'd691: color_o = 12'b000011110000;
		13'd692: color_o = 12'b000011110000;
		13'd693: color_o = 12'b000011110000;
		13'd694: color_o = 12'b000011110000;
		13'd695: color_o = 12'b000011110000;
		13'd696: color_o = 12'b000011110000;
		13'd697: color_o = 12'b000011110000;
		13'd698: color_o = 12'b000011110000;
		13'd699: color_o = 12'b000011110000;
		13'd700: color_o = 12'b000011110000;
		13'd701: color_o = 12'b000011110000;
		13'd702: color_o = 12'b000011110000;
		13'd703: color_o = 12'b000011110000;
		13'd704: color_o = 12'b000011110000;
		13'd705: color_o = 12'b000011110000;
		13'd706: color_o = 12'b000011110000;
		13'd707: color_o = 12'b000011110000;
		13'd708: color_o = 12'b000011110000;
		13'd709: color_o = 12'b000011110000;
		13'd710: color_o = 12'b000011110000;
		13'd711: color_o = 12'b000011110000;
		13'd712: color_o = 12'b000000000000;
		13'd713: color_o = 12'b000000000000;
		13'd714: color_o = 12'b100000000001;
		13'd715: color_o = 12'b000000000000;
		13'd716: color_o = 12'b100001000000;
		13'd717: color_o = 12'b100001000000;
		13'd718: color_o = 12'b100001000000;
		13'd719: color_o = 12'b100001000000;
		13'd720: color_o = 12'b000000000000;
		13'd721: color_o = 12'b100000000001;
		13'd722: color_o = 12'b100000000001;
		13'd723: color_o = 12'b000000000000;
		13'd724: color_o = 12'b000000000000;
		13'd725: color_o = 12'b000000000000;
		13'd726: color_o = 12'b000000000000;
		13'd727: color_o = 12'b000000000000;
		13'd728: color_o = 12'b000000000000;
		13'd729: color_o = 12'b000000000000;
		13'd730: color_o = 12'b000000000000;
		13'd731: color_o = 12'b000000000000;
		13'd732: color_o = 12'b000000000000;
		13'd733: color_o = 12'b000000000000;
		13'd734: color_o = 12'b000000000000;
		13'd735: color_o = 12'b000000000000;
		13'd736: color_o = 12'b000000000000;
		13'd737: color_o = 12'b000011110000;
		13'd738: color_o = 12'b000011110000;
		13'd739: color_o = 12'b000011110000;
		13'd740: color_o = 12'b000011110000;
		13'd741: color_o = 12'b000011110000;
		13'd742: color_o = 12'b000011110000;
		13'd743: color_o = 12'b000011110000;
		13'd744: color_o = 12'b000011110000;
		13'd745: color_o = 12'b000011110000;
		13'd746: color_o = 12'b000011110000;
		13'd747: color_o = 12'b000011110000;
		13'd748: color_o = 12'b000011110000;
		13'd749: color_o = 12'b000011110000;
		13'd750: color_o = 12'b000011110000;
		13'd751: color_o = 12'b000011110000;
		13'd752: color_o = 12'b000011110000;
		13'd753: color_o = 12'b000011110000;
		13'd754: color_o = 12'b000011110000;
		13'd755: color_o = 12'b000011110000;
		13'd756: color_o = 12'b000011110000;
		13'd757: color_o = 12'b000011110000;
		13'd758: color_o = 12'b000011110000;
		13'd759: color_o = 12'b000011110000;
		13'd760: color_o = 12'b000011110000;
		13'd761: color_o = 12'b000011110000;
		13'd762: color_o = 12'b000011110000;
		13'd763: color_o = 12'b000011110000;
		13'd764: color_o = 12'b000011110000;
		13'd765: color_o = 12'b000011110000;
		13'd766: color_o = 12'b000011110000;
		13'd767: color_o = 12'b000011110000;
		13'd768: color_o = 12'b000011110000;
		13'd769: color_o = 12'b000011110000;
		13'd770: color_o = 12'b000011110000;
		13'd771: color_o = 12'b000011110000;
		13'd772: color_o = 12'b000011110000;
		13'd773: color_o = 12'b000011110000;
		13'd774: color_o = 12'b000011110000;
		13'd775: color_o = 12'b000011110000;
		13'd776: color_o = 12'b000000000000;
		13'd777: color_o = 12'b000000000000;
		13'd778: color_o = 12'b100000000001;
		13'd779: color_o = 12'b000000000000;
		13'd780: color_o = 12'b100001000000;
		13'd781: color_o = 12'b100001000000;
		13'd782: color_o = 12'b100001000000;
		13'd783: color_o = 12'b100001000000;
		13'd784: color_o = 12'b000000000000;
		13'd785: color_o = 12'b100000000001;
		13'd786: color_o = 12'b100000000001;
		13'd787: color_o = 12'b000000000000;
		13'd788: color_o = 12'b000000000000;
		13'd789: color_o = 12'b000000000000;
		13'd790: color_o = 12'b000000000000;
		13'd791: color_o = 12'b000000000000;
		13'd792: color_o = 12'b000000000000;
		13'd793: color_o = 12'b000000000000;
		13'd794: color_o = 12'b110011001100;
		13'd795: color_o = 12'b110011001100;
		13'd796: color_o = 12'b110011001100;
		13'd797: color_o = 12'b000000000000;
		13'd798: color_o = 12'b000000000000;
		13'd799: color_o = 12'b000000000000;
		13'd800: color_o = 12'b000000000000;
		13'd801: color_o = 12'b000011110000;
		13'd802: color_o = 12'b000011110000;
		13'd803: color_o = 12'b000011110000;
		13'd804: color_o = 12'b000011110000;
		13'd805: color_o = 12'b000011110000;
		13'd806: color_o = 12'b000011110000;
		13'd807: color_o = 12'b000011110000;
		13'd808: color_o = 12'b000011110000;
		13'd809: color_o = 12'b000011110000;
		13'd810: color_o = 12'b000011110000;
		13'd811: color_o = 12'b000011110000;
		13'd812: color_o = 12'b000011110000;
		13'd813: color_o = 12'b000011110000;
		13'd814: color_o = 12'b000011110000;
		13'd815: color_o = 12'b000011110000;
		13'd816: color_o = 12'b000011110000;
		13'd817: color_o = 12'b000011110000;
		13'd818: color_o = 12'b000011110000;
		13'd819: color_o = 12'b000011110000;
		13'd820: color_o = 12'b000011110000;
		13'd821: color_o = 12'b000011110000;
		13'd822: color_o = 12'b000011110000;
		13'd823: color_o = 12'b000011110000;
		13'd824: color_o = 12'b000011110000;
		13'd825: color_o = 12'b000011110000;
		13'd826: color_o = 12'b000011110000;
		13'd827: color_o = 12'b000011110000;
		13'd828: color_o = 12'b000011110000;
		13'd829: color_o = 12'b000011110000;
		13'd830: color_o = 12'b000011110000;
		13'd831: color_o = 12'b000011110000;
		13'd832: color_o = 12'b000011110000;
		13'd833: color_o = 12'b000011110000;
		13'd834: color_o = 12'b000011110000;
		13'd835: color_o = 12'b000011110000;
		13'd836: color_o = 12'b000011110000;
		13'd837: color_o = 12'b000011110000;
		13'd838: color_o = 12'b000011110000;
		13'd839: color_o = 12'b000011110000;
		13'd840: color_o = 12'b000000000000;
		13'd841: color_o = 12'b100000000001;
		13'd842: color_o = 12'b100000000001;
		13'd843: color_o = 12'b000000000000;
		13'd844: color_o = 12'b100001000000;
		13'd845: color_o = 12'b100001000000;
		13'd846: color_o = 12'b100001000000;
		13'd847: color_o = 12'b100001000000;
		13'd848: color_o = 12'b000000000000;
		13'd849: color_o = 12'b100000000001;
		13'd850: color_o = 12'b000000000000;
		13'd851: color_o = 12'b000000000000;
		13'd852: color_o = 12'b000000000000;
		13'd853: color_o = 12'b000000000000;
		13'd854: color_o = 12'b000000000000;
		13'd855: color_o = 12'b000000000000;
		13'd856: color_o = 12'b000000000000;
		13'd857: color_o = 12'b000000000000;
		13'd858: color_o = 12'b110011001100;
		13'd859: color_o = 12'b110011001100;
		13'd860: color_o = 12'b110011001100;
		13'd861: color_o = 12'b000000000000;
		13'd862: color_o = 12'b000000000000;
		13'd863: color_o = 12'b000000000000;
		13'd864: color_o = 12'b000000000000;
		13'd865: color_o = 12'b000011110000;
		13'd866: color_o = 12'b000011110000;
		13'd867: color_o = 12'b000011110000;
		13'd868: color_o = 12'b000011110000;
		13'd869: color_o = 12'b000011110000;
		13'd870: color_o = 12'b000011110000;
		13'd871: color_o = 12'b000011110000;
		13'd872: color_o = 12'b000011110000;
		13'd873: color_o = 12'b000011110000;
		13'd874: color_o = 12'b000011110000;
		13'd875: color_o = 12'b000011110000;
		13'd876: color_o = 12'b000011110000;
		13'd877: color_o = 12'b000011110000;
		13'd878: color_o = 12'b000011110000;
		13'd879: color_o = 12'b000011110000;
		13'd880: color_o = 12'b000011110000;
		13'd881: color_o = 12'b000011110000;
		13'd882: color_o = 12'b000011110000;
		13'd883: color_o = 12'b000011110000;
		13'd884: color_o = 12'b000011110000;
		13'd885: color_o = 12'b000011110000;
		13'd886: color_o = 12'b000011110000;
		13'd887: color_o = 12'b000011110000;
		13'd888: color_o = 12'b000011110000;
		13'd889: color_o = 12'b000011110000;
		13'd890: color_o = 12'b000011110000;
		13'd891: color_o = 12'b000011110000;
		13'd892: color_o = 12'b000011110000;
		13'd893: color_o = 12'b000011110000;
		13'd894: color_o = 12'b000011110000;
		13'd895: color_o = 12'b000011110000;
		13'd896: color_o = 12'b000011110000;
		13'd897: color_o = 12'b000011110000;
		13'd898: color_o = 12'b000011110000;
		13'd899: color_o = 12'b000011110000;
		13'd900: color_o = 12'b000011110000;
		13'd901: color_o = 12'b000011110000;
		13'd902: color_o = 12'b000011110000;
		13'd903: color_o = 12'b000011110000;
		13'd904: color_o = 12'b000000000000;
		13'd905: color_o = 12'b100000000001;
		13'd906: color_o = 12'b100000000001;
		13'd907: color_o = 12'b000000000000;
		13'd908: color_o = 12'b000000000000;
		13'd909: color_o = 12'b000000000000;
		13'd910: color_o = 12'b100001000000;
		13'd911: color_o = 12'b100001000000;
		13'd912: color_o = 12'b000000000000;
		13'd913: color_o = 12'b100000000001;
		13'd914: color_o = 12'b100000000001;
		13'd915: color_o = 12'b000000000000;
		13'd916: color_o = 12'b000000000000;
		13'd917: color_o = 12'b000000000000;
		13'd918: color_o = 12'b000000000000;
		13'd919: color_o = 12'b000000000000;
		13'd920: color_o = 12'b000000000000;
		13'd921: color_o = 12'b000000000000;
		13'd922: color_o = 12'b000000000000;
		13'd923: color_o = 12'b000000000000;
		13'd924: color_o = 12'b110011001100;
		13'd925: color_o = 12'b000000000000;
		13'd926: color_o = 12'b000000000000;
		13'd927: color_o = 12'b000000000000;
		13'd928: color_o = 12'b000000000000;
		13'd929: color_o = 12'b000011110000;
		13'd930: color_o = 12'b000011110000;
		13'd931: color_o = 12'b000011110000;
		13'd932: color_o = 12'b000011110000;
		13'd933: color_o = 12'b000011110000;
		13'd934: color_o = 12'b000011110000;
		13'd935: color_o = 12'b000011110000;
		13'd936: color_o = 12'b000011110000;
		13'd937: color_o = 12'b000011110000;
		13'd938: color_o = 12'b000011110000;
		13'd939: color_o = 12'b000011110000;
		13'd940: color_o = 12'b000011110000;
		13'd941: color_o = 12'b000011110000;
		13'd942: color_o = 12'b000011110000;
		13'd943: color_o = 12'b000011110000;
		13'd944: color_o = 12'b000011110000;
		13'd945: color_o = 12'b000011110000;
		13'd946: color_o = 12'b000011110000;
		13'd947: color_o = 12'b000011110000;
		13'd948: color_o = 12'b000011110000;
		13'd949: color_o = 12'b000011110000;
		13'd950: color_o = 12'b000011110000;
		13'd951: color_o = 12'b000011110000;
		13'd952: color_o = 12'b000011110000;
		13'd953: color_o = 12'b000011110000;
		13'd954: color_o = 12'b000011110000;
		13'd955: color_o = 12'b000011110000;
		13'd956: color_o = 12'b000011110000;
		13'd957: color_o = 12'b000011110000;
		13'd958: color_o = 12'b000011110000;
		13'd959: color_o = 12'b000011110000;
		13'd960: color_o = 12'b000011110000;
		13'd961: color_o = 12'b000011110000;
		13'd962: color_o = 12'b000011110000;
		13'd963: color_o = 12'b000011110000;
		13'd964: color_o = 12'b000011110000;
		13'd965: color_o = 12'b000011110000;
		13'd966: color_o = 12'b000011110000;
		13'd967: color_o = 12'b000011110000;
		13'd968: color_o = 12'b100000000001;
		13'd969: color_o = 12'b100000000001;
		13'd970: color_o = 12'b100000000001;
		13'd971: color_o = 12'b100000000001;
		13'd972: color_o = 12'b000000000000;
		13'd973: color_o = 12'b000000000000;
		13'd974: color_o = 12'b000000000000;
		13'd975: color_o = 12'b000000000000;
		13'd976: color_o = 12'b000000000000;
		13'd977: color_o = 12'b000000000000;
		13'd978: color_o = 12'b100000000001;
		13'd979: color_o = 12'b100000000001;
		13'd980: color_o = 12'b000000000000;
		13'd981: color_o = 12'b000000000000;
		13'd982: color_o = 12'b000000000000;
		13'd983: color_o = 12'b000000000000;
		13'd984: color_o = 12'b000000000000;
		13'd985: color_o = 12'b000000000000;
		13'd986: color_o = 12'b000000000000;
		13'd987: color_o = 12'b000000000000;
		13'd988: color_o = 12'b000000000000;
		13'd989: color_o = 12'b000000000000;
		13'd990: color_o = 12'b000000000000;
		13'd991: color_o = 12'b000000000000;
		13'd992: color_o = 12'b000011110000;
		13'd993: color_o = 12'b000011110000;
		13'd994: color_o = 12'b000011110000;
		13'd995: color_o = 12'b000011110000;
		13'd996: color_o = 12'b000011110000;
		13'd997: color_o = 12'b000011110000;
		13'd998: color_o = 12'b000011110000;
		13'd999: color_o = 12'b000011110000;
		13'd1000: color_o = 12'b000011110000;
		13'd1001: color_o = 12'b000011110000;
		13'd1002: color_o = 12'b000011110000;
		13'd1003: color_o = 12'b000011110000;
		13'd1004: color_o = 12'b000011110000;
		13'd1005: color_o = 12'b000011110000;
		13'd1006: color_o = 12'b000011110000;
		13'd1007: color_o = 12'b000011110000;
		13'd1008: color_o = 12'b000011110000;
		13'd1009: color_o = 12'b000011110000;
		13'd1010: color_o = 12'b000011110000;
		13'd1011: color_o = 12'b000011110000;
		13'd1012: color_o = 12'b000011110000;
		13'd1013: color_o = 12'b000011110000;
		13'd1014: color_o = 12'b000011110000;
		13'd1015: color_o = 12'b000011110000;
		13'd1016: color_o = 12'b000011110000;
		13'd1017: color_o = 12'b000011110000;
		13'd1018: color_o = 12'b000011110000;
		13'd1019: color_o = 12'b000011110000;
		13'd1020: color_o = 12'b000011110000;
		13'd1021: color_o = 12'b000011110000;
		13'd1022: color_o = 12'b000011110000;
		13'd1023: color_o = 12'b000011110000;
		13'd1024: color_o = 12'b000011110000;
		13'd1025: color_o = 12'b000011110000;
		13'd1026: color_o = 12'b000011110000;
		13'd1027: color_o = 12'b000011110000;
		13'd1028: color_o = 12'b000011110000;
		13'd1029: color_o = 12'b000011110000;
		13'd1030: color_o = 12'b000011110000;
		13'd1031: color_o = 12'b000011110000;
		13'd1032: color_o = 12'b100000000001;
		13'd1033: color_o = 12'b100000000001;
		13'd1034: color_o = 12'b000000000000;
		13'd1035: color_o = 12'b000000000000;
		13'd1036: color_o = 12'b111000010010;
		13'd1037: color_o = 12'b111000010010;
		13'd1038: color_o = 12'b000000000000;
		13'd1039: color_o = 12'b000000000000;
		13'd1040: color_o = 12'b000000000000;
		13'd1041: color_o = 12'b000000000000;
		13'd1042: color_o = 12'b000000000000;
		13'd1043: color_o = 12'b000000000000;
		13'd1044: color_o = 12'b100000000001;
		13'd1045: color_o = 12'b100000000001;
		13'd1046: color_o = 12'b100000000001;
		13'd1047: color_o = 12'b100000000001;
		13'd1048: color_o = 12'b100000000001;
		13'd1049: color_o = 12'b100000000001;
		13'd1050: color_o = 12'b100000000001;
		13'd1051: color_o = 12'b100000000001;
		13'd1052: color_o = 12'b100000000001;
		13'd1053: color_o = 12'b100000000001;
		13'd1054: color_o = 12'b100000000001;
		13'd1055: color_o = 12'b100000000001;
		13'd1056: color_o = 12'b000011110000;
		13'd1057: color_o = 12'b000011110000;
		13'd1058: color_o = 12'b000011110000;
		13'd1059: color_o = 12'b000011110000;
		13'd1060: color_o = 12'b000011110000;
		13'd1061: color_o = 12'b000011110000;
		13'd1062: color_o = 12'b000011110000;
		13'd1063: color_o = 12'b000011110000;
		13'd1064: color_o = 12'b000011110000;
		13'd1065: color_o = 12'b000011110000;
		13'd1066: color_o = 12'b000011110000;
		13'd1067: color_o = 12'b000011110000;
		13'd1068: color_o = 12'b000011110000;
		13'd1069: color_o = 12'b000011110000;
		13'd1070: color_o = 12'b000011110000;
		13'd1071: color_o = 12'b000011110000;
		13'd1072: color_o = 12'b000011110000;
		13'd1073: color_o = 12'b000011110000;
		13'd1074: color_o = 12'b000011110000;
		13'd1075: color_o = 12'b000011110000;
		13'd1076: color_o = 12'b000011110000;
		13'd1077: color_o = 12'b000011110000;
		13'd1078: color_o = 12'b000011110000;
		13'd1079: color_o = 12'b000011110000;
		13'd1080: color_o = 12'b000011110000;
		13'd1081: color_o = 12'b000011110000;
		13'd1082: color_o = 12'b000011110000;
		13'd1083: color_o = 12'b000011110000;
		13'd1084: color_o = 12'b000011110000;
		13'd1085: color_o = 12'b000011110000;
		13'd1086: color_o = 12'b000011110000;
		13'd1087: color_o = 12'b000011110000;
		13'd1088: color_o = 12'b000011110000;
		13'd1089: color_o = 12'b000011110000;
		13'd1090: color_o = 12'b000011110000;
		13'd1091: color_o = 12'b000011110000;
		13'd1092: color_o = 12'b000011110000;
		13'd1093: color_o = 12'b000011110000;
		13'd1094: color_o = 12'b000011110000;
		13'd1095: color_o = 12'b000000000000;
		13'd1096: color_o = 12'b000000000000;
		13'd1097: color_o = 12'b100000000001;
		13'd1098: color_o = 12'b000000000000;
		13'd1099: color_o = 12'b111000010010;
		13'd1100: color_o = 12'b111000010010;
		13'd1101: color_o = 12'b000000000000;
		13'd1102: color_o = 12'b000000000000;
		13'd1103: color_o = 12'b100000000001;
		13'd1104: color_o = 12'b000000000000;
		13'd1105: color_o = 12'b111000010010;
		13'd1106: color_o = 12'b111000010010;
		13'd1107: color_o = 12'b000000000000;
		13'd1108: color_o = 12'b000000000000;
		13'd1109: color_o = 12'b000000000000;
		13'd1110: color_o = 12'b000000000000;
		13'd1111: color_o = 12'b000000000000;
		13'd1112: color_o = 12'b000000000000;
		13'd1113: color_o = 12'b000000000000;
		13'd1114: color_o = 12'b000000000000;
		13'd1115: color_o = 12'b000000000000;
		13'd1116: color_o = 12'b000000000000;
		13'd1117: color_o = 12'b100000000001;
		13'd1118: color_o = 12'b100000000001;
		13'd1119: color_o = 12'b100000000001;
		13'd1120: color_o = 12'b100000000001;
		13'd1121: color_o = 12'b000011110000;
		13'd1122: color_o = 12'b000011110000;
		13'd1123: color_o = 12'b000011110000;
		13'd1124: color_o = 12'b000011110000;
		13'd1125: color_o = 12'b000011110000;
		13'd1126: color_o = 12'b000011110000;
		13'd1127: color_o = 12'b000011110000;
		13'd1128: color_o = 12'b000011110000;
		13'd1129: color_o = 12'b000011110000;
		13'd1130: color_o = 12'b000011110000;
		13'd1131: color_o = 12'b000011110000;
		13'd1132: color_o = 12'b000011110000;
		13'd1133: color_o = 12'b000011110000;
		13'd1134: color_o = 12'b000011110000;
		13'd1135: color_o = 12'b000011110000;
		13'd1136: color_o = 12'b000011110000;
		13'd1137: color_o = 12'b000011110000;
		13'd1138: color_o = 12'b000011110000;
		13'd1139: color_o = 12'b000011110000;
		13'd1140: color_o = 12'b000011110000;
		13'd1141: color_o = 12'b000011110000;
		13'd1142: color_o = 12'b000011110000;
		13'd1143: color_o = 12'b000011110000;
		13'd1144: color_o = 12'b000011110000;
		13'd1145: color_o = 12'b000011110000;
		13'd1146: color_o = 12'b000011110000;
		13'd1147: color_o = 12'b000011110000;
		13'd1148: color_o = 12'b000011110000;
		13'd1149: color_o = 12'b000011110000;
		13'd1150: color_o = 12'b000011110000;
		13'd1151: color_o = 12'b000011110000;
		13'd1152: color_o = 12'b000011110000;
		13'd1153: color_o = 12'b000011110000;
		13'd1154: color_o = 12'b000011110000;
		13'd1155: color_o = 12'b000011110000;
		13'd1156: color_o = 12'b000011110000;
		13'd1157: color_o = 12'b000011110000;
		13'd1158: color_o = 12'b000000000000;
		13'd1159: color_o = 12'b000000000000;
		13'd1160: color_o = 12'b000000000000;
		13'd1161: color_o = 12'b000000000000;
		13'd1162: color_o = 12'b111000010010;
		13'd1163: color_o = 12'b111000010010;
		13'd1164: color_o = 12'b000000000000;
		13'd1165: color_o = 12'b000000000000;
		13'd1166: color_o = 12'b100000000001;
		13'd1167: color_o = 12'b100000000001;
		13'd1168: color_o = 12'b000000000000;
		13'd1169: color_o = 12'b111000010010;
		13'd1170: color_o = 12'b111000010010;
		13'd1171: color_o = 12'b000000000000;
		13'd1172: color_o = 12'b000000000000;
		13'd1173: color_o = 12'b100000000001;
		13'd1174: color_o = 12'b100000000001;
		13'd1175: color_o = 12'b100000000001;
		13'd1176: color_o = 12'b000000000000;
		13'd1177: color_o = 12'b111000010010;
		13'd1178: color_o = 12'b111000010010;
		13'd1179: color_o = 12'b000000000000;
		13'd1180: color_o = 12'b000000000000;
		13'd1181: color_o = 12'b100000000001;
		13'd1182: color_o = 12'b100000000001;
		13'd1183: color_o = 12'b100000000001;
		13'd1184: color_o = 12'b100000000001;
		13'd1185: color_o = 12'b000011110000;
		13'd1186: color_o = 12'b000011110000;
		13'd1187: color_o = 12'b000011110000;
		13'd1188: color_o = 12'b000011110000;
		13'd1189: color_o = 12'b000011110000;
		13'd1190: color_o = 12'b000011110000;
		13'd1191: color_o = 12'b000011110000;
		13'd1192: color_o = 12'b000011110000;
		13'd1193: color_o = 12'b000011110000;
		13'd1194: color_o = 12'b000011110000;
		13'd1195: color_o = 12'b000011110000;
		13'd1196: color_o = 12'b000011110000;
		13'd1197: color_o = 12'b000011110000;
		13'd1198: color_o = 12'b000011110000;
		13'd1199: color_o = 12'b000011110000;
		13'd1200: color_o = 12'b000011110000;
		13'd1201: color_o = 12'b000011110000;
		13'd1202: color_o = 12'b000011110000;
		13'd1203: color_o = 12'b000011110000;
		13'd1204: color_o = 12'b000011110000;
		13'd1205: color_o = 12'b000011110000;
		13'd1206: color_o = 12'b000011110000;
		13'd1207: color_o = 12'b000011110000;
		13'd1208: color_o = 12'b000011110000;
		13'd1209: color_o = 12'b000011110000;
		13'd1210: color_o = 12'b000011110000;
		13'd1211: color_o = 12'b000011110000;
		13'd1212: color_o = 12'b000011110000;
		13'd1213: color_o = 12'b000011110000;
		13'd1214: color_o = 12'b000011110000;
		13'd1215: color_o = 12'b000011110000;
		13'd1216: color_o = 12'b000011110000;
		13'd1217: color_o = 12'b000011110000;
		13'd1218: color_o = 12'b000011110000;
		13'd1219: color_o = 12'b000011110000;
		13'd1220: color_o = 12'b000011110000;
		13'd1221: color_o = 12'b000000000000;
		13'd1222: color_o = 12'b000000000000;
		13'd1223: color_o = 12'b000000000000;
		13'd1224: color_o = 12'b000000000000;
		13'd1225: color_o = 12'b100000000000;
		13'd1226: color_o = 12'b100000000000;
		13'd1227: color_o = 12'b100000000001;
		13'd1228: color_o = 12'b000000000000;
		13'd1229: color_o = 12'b100000000001;
		13'd1230: color_o = 12'b100000000001;
		13'd1231: color_o = 12'b000000000000;
		13'd1232: color_o = 12'b000000000000;
		13'd1233: color_o = 12'b000000000000;
		13'd1234: color_o = 12'b000000000000;
		13'd1235: color_o = 12'b000000000000;
		13'd1236: color_o = 12'b000000000000;
		13'd1237: color_o = 12'b000000000000;
		13'd1238: color_o = 12'b000000000000;
		13'd1239: color_o = 12'b000000000000;
		13'd1240: color_o = 12'b111000010010;
		13'd1241: color_o = 12'b111000010010;
		13'd1242: color_o = 12'b111000010010;
		13'd1243: color_o = 12'b000000000000;
		13'd1244: color_o = 12'b100000000001;
		13'd1245: color_o = 12'b100000000001;
		13'd1246: color_o = 12'b100000000001;
		13'd1247: color_o = 12'b100000000001;
		13'd1248: color_o = 12'b000000000000;
		13'd1249: color_o = 12'b000011110000;
		13'd1250: color_o = 12'b000011110000;
		13'd1251: color_o = 12'b000011110000;
		13'd1252: color_o = 12'b000011110000;
		13'd1253: color_o = 12'b000011110000;
		13'd1254: color_o = 12'b000011110000;
		13'd1255: color_o = 12'b000011110000;
		13'd1256: color_o = 12'b000011110000;
		13'd1257: color_o = 12'b000011110000;
		13'd1258: color_o = 12'b000011110000;
		13'd1259: color_o = 12'b000011110000;
		13'd1260: color_o = 12'b000011110000;
		13'd1261: color_o = 12'b000011110000;
		13'd1262: color_o = 12'b000011110000;
		13'd1263: color_o = 12'b000011110000;
		13'd1264: color_o = 12'b000011110000;
		13'd1265: color_o = 12'b000011110000;
		13'd1266: color_o = 12'b000011110000;
		13'd1267: color_o = 12'b000011110000;
		13'd1268: color_o = 12'b000011110000;
		13'd1269: color_o = 12'b000011110000;
		13'd1270: color_o = 12'b000011110000;
		13'd1271: color_o = 12'b000011110000;
		13'd1272: color_o = 12'b000011110000;
		13'd1273: color_o = 12'b000011110000;
		13'd1274: color_o = 12'b000011110000;
		13'd1275: color_o = 12'b000011110000;
		13'd1276: color_o = 12'b000011110000;
		13'd1277: color_o = 12'b000011110000;
		13'd1278: color_o = 12'b000011110000;
		13'd1279: color_o = 12'b000011110000;
		13'd1280: color_o = 12'b000011110000;
		13'd1281: color_o = 12'b000011110000;
		13'd1282: color_o = 12'b000011110000;
		13'd1283: color_o = 12'b000011110000;
		13'd1284: color_o = 12'b000011110000;
		13'd1285: color_o = 12'b000000000000;
		13'd1286: color_o = 12'b100001000000;
		13'd1287: color_o = 12'b000000000000;
		13'd1288: color_o = 12'b000000000000;
		13'd1289: color_o = 12'b100000000001;
		13'd1290: color_o = 12'b100000000001;
		13'd1291: color_o = 12'b100000000000;
		13'd1292: color_o = 12'b000000000000;
		13'd1293: color_o = 12'b000000000000;
		13'd1294: color_o = 12'b000000000000;
		13'd1295: color_o = 12'b000000000000;
		13'd1296: color_o = 12'b100000000000;
		13'd1297: color_o = 12'b100000000000;
		13'd1298: color_o = 12'b100000000000;
		13'd1299: color_o = 12'b000000000000;
		13'd1300: color_o = 12'b000000000000;
		13'd1301: color_o = 12'b000000000000;
		13'd1302: color_o = 12'b000000000000;
		13'd1303: color_o = 12'b000000000000;
		13'd1304: color_o = 12'b000000000000;
		13'd1305: color_o = 12'b111000010010;
		13'd1306: color_o = 12'b111000010010;
		13'd1307: color_o = 12'b000000000000;
		13'd1308: color_o = 12'b000000000000;
		13'd1309: color_o = 12'b000000000000;
		13'd1310: color_o = 12'b000000000000;
		13'd1311: color_o = 12'b000000000000;
		13'd1312: color_o = 12'b000000000000;
		13'd1313: color_o = 12'b000011110000;
		13'd1314: color_o = 12'b000011110000;
		13'd1315: color_o = 12'b000011110000;
		13'd1316: color_o = 12'b000011110000;
		13'd1317: color_o = 12'b000011110000;
		13'd1318: color_o = 12'b000011110000;
		13'd1319: color_o = 12'b000011110000;
		13'd1320: color_o = 12'b000011110000;
		13'd1321: color_o = 12'b000011110000;
		13'd1322: color_o = 12'b000011110000;
		13'd1323: color_o = 12'b000011110000;
		13'd1324: color_o = 12'b000011110000;
		13'd1325: color_o = 12'b000011110000;
		13'd1326: color_o = 12'b000011110000;
		13'd1327: color_o = 12'b000011110000;
		13'd1328: color_o = 12'b000011110000;
		13'd1329: color_o = 12'b000011110000;
		13'd1330: color_o = 12'b000011110000;
		13'd1331: color_o = 12'b000011110000;
		13'd1332: color_o = 12'b000011110000;
		13'd1333: color_o = 12'b000011110000;
		13'd1334: color_o = 12'b000011110000;
		13'd1335: color_o = 12'b000011110000;
		13'd1336: color_o = 12'b000011110000;
		13'd1337: color_o = 12'b000011110000;
		13'd1338: color_o = 12'b000011110000;
		13'd1339: color_o = 12'b000011110000;
		13'd1340: color_o = 12'b000011110000;
		13'd1341: color_o = 12'b000011110000;
		13'd1342: color_o = 12'b000011110000;
		13'd1343: color_o = 12'b000011110000;
		13'd1344: color_o = 12'b000011110000;
		13'd1345: color_o = 12'b000011110000;
		13'd1346: color_o = 12'b000011110000;
		13'd1347: color_o = 12'b000011110000;
		13'd1348: color_o = 12'b000000000000;
		13'd1349: color_o = 12'b000000000000;
		13'd1350: color_o = 12'b100001000000;
		13'd1351: color_o = 12'b000000000000;
		13'd1352: color_o = 12'b000000000000;
		13'd1353: color_o = 12'b100000000001;
		13'd1354: color_o = 12'b100000000001;
		13'd1355: color_o = 12'b100000000000;
		13'd1356: color_o = 12'b100000000000;
		13'd1357: color_o = 12'b000000000000;
		13'd1358: color_o = 12'b000000000000;
		13'd1359: color_o = 12'b100000000000;
		13'd1360: color_o = 12'b100000000000;
		13'd1361: color_o = 12'b100000000000;
		13'd1362: color_o = 12'b100000000000;
		13'd1363: color_o = 12'b100000000000;
		13'd1364: color_o = 12'b100000000000;
		13'd1365: color_o = 12'b100000000000;
		13'd1366: color_o = 12'b000000000000;
		13'd1367: color_o = 12'b000000000000;
		13'd1368: color_o = 12'b000000000000;
		13'd1369: color_o = 12'b000000000000;
		13'd1370: color_o = 12'b000000000000;
		13'd1371: color_o = 12'b000000000000;
		13'd1372: color_o = 12'b000000000000;
		13'd1373: color_o = 12'b000011110000;
		13'd1374: color_o = 12'b000011110000;
		13'd1375: color_o = 12'b000011110000;
		13'd1376: color_o = 12'b000011110000;
		13'd1377: color_o = 12'b000011110000;
		13'd1378: color_o = 12'b000011110000;
		13'd1379: color_o = 12'b000011110000;
		13'd1380: color_o = 12'b000011110000;
		13'd1381: color_o = 12'b000011110000;
		13'd1382: color_o = 12'b000011110000;
		13'd1383: color_o = 12'b000011110000;
		13'd1384: color_o = 12'b000011110000;
		13'd1385: color_o = 12'b000011110000;
		13'd1386: color_o = 12'b000011110000;
		13'd1387: color_o = 12'b000011110000;
		13'd1388: color_o = 12'b000011110000;
		13'd1389: color_o = 12'b000011110000;
		13'd1390: color_o = 12'b000011110000;
		13'd1391: color_o = 12'b000011110000;
		13'd1392: color_o = 12'b000011110000;
		13'd1393: color_o = 12'b000011110000;
		13'd1394: color_o = 12'b000011110000;
		13'd1395: color_o = 12'b000011110000;
		13'd1396: color_o = 12'b000011110000;
		13'd1397: color_o = 12'b000011110000;
		13'd1398: color_o = 12'b000011110000;
		13'd1399: color_o = 12'b000011110000;
		13'd1400: color_o = 12'b000011110000;
		13'd1401: color_o = 12'b000011110000;
		13'd1402: color_o = 12'b000011110000;
		13'd1403: color_o = 12'b000011110000;
		13'd1404: color_o = 12'b000011110000;
		13'd1405: color_o = 12'b000011110000;
		13'd1406: color_o = 12'b000011110000;
		13'd1407: color_o = 12'b000011110000;
		13'd1408: color_o = 12'b000011110000;
		13'd1409: color_o = 12'b000011110000;
		13'd1410: color_o = 12'b000011110000;
		13'd1411: color_o = 12'b000011110000;
		13'd1412: color_o = 12'b000000000000;
		13'd1413: color_o = 12'b100000000001;
		13'd1414: color_o = 12'b000000000000;
		13'd1415: color_o = 12'b000000000000;
		13'd1416: color_o = 12'b000000000000;
		13'd1417: color_o = 12'b100000000001;
		13'd1418: color_o = 12'b100000000001;
		13'd1419: color_o = 12'b100000000001;
		13'd1420: color_o = 12'b100000000000;
		13'd1421: color_o = 12'b000000000000;
		13'd1422: color_o = 12'b100000000000;
		13'd1423: color_o = 12'b100000000000;
		13'd1424: color_o = 12'b000000000000;
		13'd1425: color_o = 12'b100000000000;
		13'd1426: color_o = 12'b100000000000;
		13'd1427: color_o = 12'b100000000000;
		13'd1428: color_o = 12'b100000000000;
		13'd1429: color_o = 12'b100000000000;
		13'd1430: color_o = 12'b000000000000;
		13'd1431: color_o = 12'b100000000000;
		13'd1432: color_o = 12'b000000000000;
		13'd1433: color_o = 12'b000000000000;
		13'd1434: color_o = 12'b000000000000;
		13'd1435: color_o = 12'b000000000000;
		13'd1436: color_o = 12'b000000000000;
		13'd1437: color_o = 12'b000011110000;
		13'd1438: color_o = 12'b000011110000;
		13'd1439: color_o = 12'b000011110000;
		13'd1440: color_o = 12'b000011110000;
		13'd1441: color_o = 12'b000011110000;
		13'd1442: color_o = 12'b000011110000;
		13'd1443: color_o = 12'b000011110000;
		13'd1444: color_o = 12'b000011110000;
		13'd1445: color_o = 12'b000011110000;
		13'd1446: color_o = 12'b000011110000;
		13'd1447: color_o = 12'b000011110000;
		13'd1448: color_o = 12'b000011110000;
		13'd1449: color_o = 12'b000011110000;
		13'd1450: color_o = 12'b000011110000;
		13'd1451: color_o = 12'b000011110000;
		13'd1452: color_o = 12'b000011110000;
		13'd1453: color_o = 12'b000011110000;
		13'd1454: color_o = 12'b000011110000;
		13'd1455: color_o = 12'b000011110000;
		13'd1456: color_o = 12'b000011110000;
		13'd1457: color_o = 12'b000011110000;
		13'd1458: color_o = 12'b000011110000;
		13'd1459: color_o = 12'b000011110000;
		13'd1460: color_o = 12'b000011110000;
		13'd1461: color_o = 12'b000011110000;
		13'd1462: color_o = 12'b000011110000;
		13'd1463: color_o = 12'b000011110000;
		13'd1464: color_o = 12'b000011110000;
		13'd1465: color_o = 12'b000011110000;
		13'd1466: color_o = 12'b000011110000;
		13'd1467: color_o = 12'b000011110000;
		13'd1468: color_o = 12'b000011110000;
		13'd1469: color_o = 12'b000011110000;
		13'd1470: color_o = 12'b000011110000;
		13'd1471: color_o = 12'b000011110000;
		13'd1472: color_o = 12'b000011110000;
		13'd1473: color_o = 12'b000011110000;
		13'd1474: color_o = 12'b000011110000;
		13'd1475: color_o = 12'b000011110000;
		13'd1476: color_o = 12'b000000000000;
		13'd1477: color_o = 12'b100000000001;
		13'd1478: color_o = 12'b000000000000;
		13'd1479: color_o = 12'b100000000000;
		13'd1480: color_o = 12'b000000000000;
		13'd1481: color_o = 12'b100000000001;
		13'd1482: color_o = 12'b100000000001;
		13'd1483: color_o = 12'b100000000001;
		13'd1484: color_o = 12'b100000000000;
		13'd1485: color_o = 12'b000000000000;
		13'd1486: color_o = 12'b100000000000;
		13'd1487: color_o = 12'b100000000000;
		13'd1488: color_o = 12'b000000000000;
		13'd1489: color_o = 12'b000000000000;
		13'd1490: color_o = 12'b100000000000;
		13'd1491: color_o = 12'b000000000000;
		13'd1492: color_o = 12'b000000000000;
		13'd1493: color_o = 12'b100000000000;
		13'd1494: color_o = 12'b000000000000;
		13'd1495: color_o = 12'b100000000000;
		13'd1496: color_o = 12'b000000000000;
		13'd1497: color_o = 12'b100000000000;
		13'd1498: color_o = 12'b100000000000;
		13'd1499: color_o = 12'b100000000000;
		13'd1500: color_o = 12'b000000000000;
		13'd1501: color_o = 12'b000000000000;
		13'd1502: color_o = 12'b000000000000;
		13'd1503: color_o = 12'b000000000000;
		13'd1504: color_o = 12'b000011110000;
		13'd1505: color_o = 12'b000011110000;
		13'd1506: color_o = 12'b000011110000;
		13'd1507: color_o = 12'b000011110000;
		13'd1508: color_o = 12'b000011110000;
		13'd1509: color_o = 12'b000011110000;
		13'd1510: color_o = 12'b000000000000;
		13'd1511: color_o = 12'b000000000000;
		13'd1512: color_o = 12'b000000000000;
		13'd1513: color_o = 12'b000000000000;
		13'd1514: color_o = 12'b000000000000;
		13'd1515: color_o = 12'b000000000000;
		13'd1516: color_o = 12'b000000000000;
		13'd1517: color_o = 12'b000000000000;
		13'd1518: color_o = 12'b000000000000;
		13'd1519: color_o = 12'b000000000000;
		13'd1520: color_o = 12'b000000000000;
		13'd1521: color_o = 12'b000000000000;
		13'd1522: color_o = 12'b000000000000;
		13'd1523: color_o = 12'b000000000000;
		13'd1524: color_o = 12'b000000000000;
		13'd1525: color_o = 12'b000000000000;
		13'd1526: color_o = 12'b000011110000;
		13'd1527: color_o = 12'b000011110000;
		13'd1528: color_o = 12'b000011110000;
		13'd1529: color_o = 12'b000011110000;
		13'd1530: color_o = 12'b000011110000;
		13'd1531: color_o = 12'b000011110000;
		13'd1532: color_o = 12'b000011110000;
		13'd1533: color_o = 12'b000011110000;
		13'd1534: color_o = 12'b000011110000;
		13'd1535: color_o = 12'b000011110000;
		13'd1536: color_o = 12'b000011110000;
		13'd1537: color_o = 12'b000011110000;
		13'd1538: color_o = 12'b000011110000;
		13'd1539: color_o = 12'b000000000000;
		13'd1540: color_o = 12'b000000000000;
		13'd1541: color_o = 12'b100000000001;
		13'd1542: color_o = 12'b000000000000;
		13'd1543: color_o = 12'b000000000000;
		13'd1544: color_o = 12'b000000000000;
		13'd1545: color_o = 12'b100000000001;
		13'd1546: color_o = 12'b100000000001;
		13'd1547: color_o = 12'b100000000000;
		13'd1548: color_o = 12'b100000000000;
		13'd1549: color_o = 12'b000000000000;
		13'd1550: color_o = 12'b100000000000;
		13'd1551: color_o = 12'b100000000000;
		13'd1552: color_o = 12'b100000000000;
		13'd1553: color_o = 12'b000000000000;
		13'd1554: color_o = 12'b000000000000;
		13'd1555: color_o = 12'b000000000000;
		13'd1556: color_o = 12'b000000000000;
		13'd1557: color_o = 12'b100000000000;
		13'd1558: color_o = 12'b000000000000;
		13'd1559: color_o = 12'b100000000000;
		13'd1560: color_o = 12'b000000000000;
		13'd1561: color_o = 12'b000000000000;
		13'd1562: color_o = 12'b100000000000;
		13'd1563: color_o = 12'b100000000000;
		13'd1564: color_o = 12'b100000000000;
		13'd1565: color_o = 12'b000000000000;
		13'd1566: color_o = 12'b000000000000;
		13'd1567: color_o = 12'b100000000000;
		13'd1568: color_o = 12'b100000000000;
		13'd1569: color_o = 12'b000011110000;
		13'd1570: color_o = 12'b000011110000;
		13'd1571: color_o = 12'b000011110000;
		13'd1572: color_o = 12'b000000000000;
		13'd1573: color_o = 12'b000000000000;
		13'd1574: color_o = 12'b011110011011;
		13'd1575: color_o = 12'b010001000100;
		13'd1576: color_o = 12'b010001000100;
		13'd1577: color_o = 12'b010001000100;
		13'd1578: color_o = 12'b010001000100;
		13'd1579: color_o = 12'b010001000100;
		13'd1580: color_o = 12'b010001000100;
		13'd1581: color_o = 12'b010001000100;
		13'd1582: color_o = 12'b010001000100;
		13'd1583: color_o = 12'b010001000100;
		13'd1584: color_o = 12'b010001000100;
		13'd1585: color_o = 12'b010001000100;
		13'd1586: color_o = 12'b010001000100;
		13'd1587: color_o = 12'b010001000100;
		13'd1588: color_o = 12'b010001000100;
		13'd1589: color_o = 12'b010001000100;
		13'd1590: color_o = 12'b000011110000;
		13'd1591: color_o = 12'b000011110000;
		13'd1592: color_o = 12'b000011110000;
		13'd1593: color_o = 12'b000011110000;
		13'd1594: color_o = 12'b000011110000;
		13'd1595: color_o = 12'b000011110000;
		13'd1596: color_o = 12'b000011110000;
		13'd1597: color_o = 12'b000011110000;
		13'd1598: color_o = 12'b000011110000;
		13'd1599: color_o = 12'b000011110000;
		13'd1600: color_o = 12'b000011110000;
		13'd1601: color_o = 12'b000011110000;
		13'd1602: color_o = 12'b000011110000;
		13'd1603: color_o = 12'b000000000000;
		13'd1604: color_o = 12'b100000000001;
		13'd1605: color_o = 12'b100000000001;
		13'd1606: color_o = 12'b000000000000;
		13'd1607: color_o = 12'b100000000000;
		13'd1608: color_o = 12'b000000000000;
		13'd1609: color_o = 12'b100000000001;
		13'd1610: color_o = 12'b100000000001;
		13'd1611: color_o = 12'b100000000000;
		13'd1612: color_o = 12'b100000000000;
		13'd1613: color_o = 12'b000000000000;
		13'd1614: color_o = 12'b100000000000;
		13'd1615: color_o = 12'b100000000000;
		13'd1616: color_o = 12'b100000000000;
		13'd1617: color_o = 12'b000000000000;
		13'd1618: color_o = 12'b000000000000;
		13'd1619: color_o = 12'b000000000000;
		13'd1620: color_o = 12'b000000000000;
		13'd1621: color_o = 12'b100000000000;
		13'd1622: color_o = 12'b000000000000;
		13'd1623: color_o = 12'b100000000000;
		13'd1624: color_o = 12'b000000000000;
		13'd1625: color_o = 12'b100000000000;
		13'd1626: color_o = 12'b000000000000;
		13'd1627: color_o = 12'b000000000000;
		13'd1628: color_o = 12'b000000000000;
		13'd1629: color_o = 12'b000000000000;
		13'd1630: color_o = 12'b000000000000;
		13'd1631: color_o = 12'b000000000000;
		13'd1632: color_o = 12'b000000000000;
		13'd1633: color_o = 12'b000000000000;
		13'd1634: color_o = 12'b000000000000;
		13'd1635: color_o = 12'b000000000000;
		13'd1636: color_o = 12'b011110011011;
		13'd1637: color_o = 12'b011110011011;
		13'd1638: color_o = 12'b011110011011;
		13'd1639: color_o = 12'b011101110111;
		13'd1640: color_o = 12'b011101110111;
		13'd1641: color_o = 12'b011101110111;
		13'd1642: color_o = 12'b011101110111;
		13'd1643: color_o = 12'b011101110111;
		13'd1644: color_o = 12'b011101110111;
		13'd1645: color_o = 12'b011101110111;
		13'd1646: color_o = 12'b011101110111;
		13'd1647: color_o = 12'b011101110111;
		13'd1648: color_o = 12'b011101110111;
		13'd1649: color_o = 12'b011101110111;
		13'd1650: color_o = 12'b011101110111;
		13'd1651: color_o = 12'b011101110111;
		13'd1652: color_o = 12'b011101110111;
		13'd1653: color_o = 12'b011101110111;
		13'd1654: color_o = 12'b000011110000;
		13'd1655: color_o = 12'b000011110000;
		13'd1656: color_o = 12'b000011110000;
		13'd1657: color_o = 12'b000011110000;
		13'd1658: color_o = 12'b000011110000;
		13'd1659: color_o = 12'b000011110000;
		13'd1660: color_o = 12'b000011110000;
		13'd1661: color_o = 12'b000011110000;
		13'd1662: color_o = 12'b000011110000;
		13'd1663: color_o = 12'b000011110000;
		13'd1664: color_o = 12'b000011110000;
		13'd1665: color_o = 12'b000011110000;
		13'd1666: color_o = 12'b000000000000;
		13'd1667: color_o = 12'b000000000000;
		13'd1668: color_o = 12'b100000000001;
		13'd1669: color_o = 12'b100000000001;
		13'd1670: color_o = 12'b000000000000;
		13'd1671: color_o = 12'b100000000000;
		13'd1672: color_o = 12'b000000000000;
		13'd1673: color_o = 12'b000000000000;
		13'd1674: color_o = 12'b100000000001;
		13'd1675: color_o = 12'b100000000001;
		13'd1676: color_o = 12'b100000000000;
		13'd1677: color_o = 12'b000000000000;
		13'd1678: color_o = 12'b100000000000;
		13'd1679: color_o = 12'b000000000000;
		13'd1680: color_o = 12'b000000000000;
		13'd1681: color_o = 12'b000000000000;
		13'd1682: color_o = 12'b000000000000;
		13'd1683: color_o = 12'b000000000000;
		13'd1684: color_o = 12'b000000000000;
		13'd1685: color_o = 12'b100000000000;
		13'd1686: color_o = 12'b000000000000;
		13'd1687: color_o = 12'b100000000000;
		13'd1688: color_o = 12'b000000000000;
		13'd1689: color_o = 12'b100000000000;
		13'd1690: color_o = 12'b100000000000;
		13'd1691: color_o = 12'b000000000000;
		13'd1692: color_o = 12'b010001000100;
		13'd1693: color_o = 12'b010001000100;
		13'd1694: color_o = 12'b010001000100;
		13'd1695: color_o = 12'b010001000100;
		13'd1696: color_o = 12'b010001000100;
		13'd1697: color_o = 12'b010001000100;
		13'd1698: color_o = 12'b010001000100;
		13'd1699: color_o = 12'b010001000100;
		13'd1700: color_o = 12'b010001000100;
		13'd1701: color_o = 12'b010001000100;
		13'd1702: color_o = 12'b000000000000;
		13'd1703: color_o = 12'b000000000000;
		13'd1704: color_o = 12'b000000000000;
		13'd1705: color_o = 12'b000000000000;
		13'd1706: color_o = 12'b000000000000;
		13'd1707: color_o = 12'b000000000000;
		13'd1708: color_o = 12'b000000000000;
		13'd1709: color_o = 12'b000000000000;
		13'd1710: color_o = 12'b000000000000;
		13'd1711: color_o = 12'b000000000000;
		13'd1712: color_o = 12'b000000000000;
		13'd1713: color_o = 12'b000000000000;
		13'd1714: color_o = 12'b000000000000;
		13'd1715: color_o = 12'b000000000000;
		13'd1716: color_o = 12'b000000000000;
		13'd1717: color_o = 12'b000000000000;
		13'd1718: color_o = 12'b010001000100;
		13'd1719: color_o = 12'b000011110000;
		13'd1720: color_o = 12'b000011110000;
		13'd1721: color_o = 12'b000011110000;
		13'd1722: color_o = 12'b000011110000;
		13'd1723: color_o = 12'b000011110000;
		13'd1724: color_o = 12'b000011110000;
		13'd1725: color_o = 12'b000011110000;
		13'd1726: color_o = 12'b000011110000;
		13'd1727: color_o = 12'b000011110000;
		13'd1728: color_o = 12'b000011110000;
		13'd1729: color_o = 12'b000011110000;
		13'd1730: color_o = 12'b000000000000;
		13'd1731: color_o = 12'b000000000000;
		13'd1732: color_o = 12'b100000000001;
		13'd1733: color_o = 12'b100000000001;
		13'd1734: color_o = 12'b000000000000;
		13'd1735: color_o = 12'b100000000000;
		13'd1736: color_o = 12'b100000000000;
		13'd1737: color_o = 12'b100000000000;
		13'd1738: color_o = 12'b000000000000;
		13'd1739: color_o = 12'b100000000000;
		13'd1740: color_o = 12'b100000000000;
		13'd1741: color_o = 12'b000000000000;
		13'd1742: color_o = 12'b000000000000;
		13'd1743: color_o = 12'b000000000000;
		13'd1744: color_o = 12'b100000000000;
		13'd1745: color_o = 12'b100000000000;
		13'd1746: color_o = 12'b100000000000;
		13'd1747: color_o = 12'b100000000000;
		13'd1748: color_o = 12'b100000000000;
		13'd1749: color_o = 12'b100000000000;
		13'd1750: color_o = 12'b100000000000;
		13'd1751: color_o = 12'b100000000000;
		13'd1752: color_o = 12'b000000000000;
		13'd1753: color_o = 12'b100000000000;
		13'd1754: color_o = 12'b100000000000;
		13'd1755: color_o = 12'b000000000000;
		13'd1756: color_o = 12'b011110011011;
		13'd1757: color_o = 12'b011110011011;
		13'd1758: color_o = 12'b011101110111;
		13'd1759: color_o = 12'b011101110111;
		13'd1760: color_o = 12'b011101110111;
		13'd1761: color_o = 12'b011101110111;
		13'd1762: color_o = 12'b011101110111;
		13'd1763: color_o = 12'b011101110111;
		13'd1764: color_o = 12'b011101110111;
		13'd1765: color_o = 12'b011101110111;
		13'd1766: color_o = 12'b001101000110;
		13'd1767: color_o = 12'b011110011011;
		13'd1768: color_o = 12'b011110011011;
		13'd1769: color_o = 12'b011110011011;
		13'd1770: color_o = 12'b011101110111;
		13'd1771: color_o = 12'b011101110111;
		13'd1772: color_o = 12'b011101110111;
		13'd1773: color_o = 12'b011101110111;
		13'd1774: color_o = 12'b011110011011;
		13'd1775: color_o = 12'b011110011011;
		13'd1776: color_o = 12'b011101110111;
		13'd1777: color_o = 12'b011101110111;
		13'd1778: color_o = 12'b011101110111;
		13'd1779: color_o = 12'b011101110111;
		13'd1780: color_o = 12'b011101110111;
		13'd1781: color_o = 12'b011101110111;
		13'd1782: color_o = 12'b010001000100;
		13'd1783: color_o = 12'b000011110000;
		13'd1784: color_o = 12'b000011110000;
		13'd1785: color_o = 12'b000011110000;
		13'd1786: color_o = 12'b000011110000;
		13'd1787: color_o = 12'b000011110000;
		13'd1788: color_o = 12'b000011110000;
		13'd1789: color_o = 12'b000011110000;
		13'd1790: color_o = 12'b000011110000;
		13'd1791: color_o = 12'b000011110000;
		13'd1792: color_o = 12'b000011110000;
		13'd1793: color_o = 12'b000011110000;
		13'd1794: color_o = 12'b000000000000;
		13'd1795: color_o = 12'b000000000000;
		13'd1796: color_o = 12'b100000000001;
		13'd1797: color_o = 12'b100000000001;
		13'd1798: color_o = 12'b000000000000;
		13'd1799: color_o = 12'b000000000000;
		13'd1800: color_o = 12'b100000000000;
		13'd1801: color_o = 12'b100000000000;
		13'd1802: color_o = 12'b000000000000;
		13'd1803: color_o = 12'b100000000000;
		13'd1804: color_o = 12'b000000000000;
		13'd1805: color_o = 12'b000000000000;
		13'd1806: color_o = 12'b000000000000;
		13'd1807: color_o = 12'b000000000000;
		13'd1808: color_o = 12'b000000000000;
		13'd1809: color_o = 12'b000000000000;
		13'd1810: color_o = 12'b000000000000;
		13'd1811: color_o = 12'b000000000000;
		13'd1812: color_o = 12'b100000000000;
		13'd1813: color_o = 12'b100000000000;
		13'd1814: color_o = 12'b100000000000;
		13'd1815: color_o = 12'b100000000000;
		13'd1816: color_o = 12'b100000000000;
		13'd1817: color_o = 12'b100000000000;
		13'd1818: color_o = 12'b100000000000;
		13'd1819: color_o = 12'b000000000000;
		13'd1820: color_o = 12'b100000000000;
		13'd1821: color_o = 12'b000000000000;
		13'd1822: color_o = 12'b000000000000;
		13'd1823: color_o = 12'b000000000000;
		13'd1824: color_o = 12'b000000000000;
		13'd1825: color_o = 12'b000000000000;
		13'd1826: color_o = 12'b100000000000;
		13'd1827: color_o = 12'b000000000000;
		13'd1828: color_o = 12'b000000000000;
		13'd1829: color_o = 12'b100000000001;
		13'd1830: color_o = 12'b100000000001;
		13'd1831: color_o = 12'b100000000001;
		13'd1832: color_o = 12'b011101110111;
		13'd1833: color_o = 12'b011101110111;
		13'd1834: color_o = 12'b011101110111;
		13'd1835: color_o = 12'b011110011011;
		13'd1836: color_o = 12'b011110011011;
		13'd1837: color_o = 12'b011110011011;
		13'd1838: color_o = 12'b011101110111;
		13'd1839: color_o = 12'b011101110111;
		13'd1840: color_o = 12'b011101110111;
		13'd1841: color_o = 12'b011110011011;
		13'd1842: color_o = 12'b011010001010;
		13'd1843: color_o = 12'b011110011011;
		13'd1844: color_o = 12'b011101110111;
		13'd1845: color_o = 12'b011101110111;
		13'd1846: color_o = 12'b011101110111;
		13'd1847: color_o = 12'b010001000100;
		13'd1848: color_o = 12'b000011110000;
		13'd1849: color_o = 12'b000011110000;
		13'd1850: color_o = 12'b000011110000;
		13'd1851: color_o = 12'b000011110000;
		13'd1852: color_o = 12'b000011110000;
		13'd1853: color_o = 12'b000011110000;
		13'd1854: color_o = 12'b000011110000;
		13'd1855: color_o = 12'b000011110000;
		13'd1856: color_o = 12'b000011110000;
		13'd1857: color_o = 12'b000011110000;
		13'd1858: color_o = 12'b000000000000;
		13'd1859: color_o = 12'b000000000000;
		13'd1860: color_o = 12'b100000000001;
		13'd1861: color_o = 12'b100000000001;
		13'd1862: color_o = 12'b100000000001;
		13'd1863: color_o = 12'b000000000000;
		13'd1864: color_o = 12'b100000000000;
		13'd1865: color_o = 12'b000000000000;
		13'd1866: color_o = 12'b000000000000;
		13'd1867: color_o = 12'b100000000000;
		13'd1868: color_o = 12'b100000000000;
		13'd1869: color_o = 12'b000000000000;
		13'd1870: color_o = 12'b000000000000;
		13'd1871: color_o = 12'b000000000000;
		13'd1872: color_o = 12'b100000000001;
		13'd1873: color_o = 12'b100000000001;
		13'd1874: color_o = 12'b100000000001;
		13'd1875: color_o = 12'b100000000001;
		13'd1876: color_o = 12'b100000000000;
		13'd1877: color_o = 12'b100000000001;
		13'd1878: color_o = 12'b100000000001;
		13'd1879: color_o = 12'b100000000001;
		13'd1880: color_o = 12'b100000000000;
		13'd1881: color_o = 12'b100000000000;
		13'd1882: color_o = 12'b000000000000;
		13'd1883: color_o = 12'b000000000000;
		13'd1884: color_o = 12'b100000000000;
		13'd1885: color_o = 12'b100000000000;
		13'd1886: color_o = 12'b100000000000;
		13'd1887: color_o = 12'b100000000000;
		13'd1888: color_o = 12'b100000000000;
		13'd1889: color_o = 12'b100000000000;
		13'd1890: color_o = 12'b100000000000;
		13'd1891: color_o = 12'b100000000000;
		13'd1892: color_o = 12'b000000000000;
		13'd1893: color_o = 12'b000000000000;
		13'd1894: color_o = 12'b100000000001;
		13'd1895: color_o = 12'b000000000000;
		13'd1896: color_o = 12'b000000000000;
		13'd1897: color_o = 12'b000000000000;
		13'd1898: color_o = 12'b000000000000;
		13'd1899: color_o = 12'b000000000000;
		13'd1900: color_o = 12'b000000000000;
		13'd1901: color_o = 12'b000000000000;
		13'd1902: color_o = 12'b000000000000;
		13'd1903: color_o = 12'b000000000000;
		13'd1904: color_o = 12'b000000000000;
		13'd1905: color_o = 12'b000000000000;
		13'd1906: color_o = 12'b000000000000;
		13'd1907: color_o = 12'b000000000000;
		13'd1908: color_o = 12'b011110011011;
		13'd1909: color_o = 12'b011101110111;
		13'd1910: color_o = 12'b011101110111;
		13'd1911: color_o = 12'b011101110111;
		13'd1912: color_o = 12'b000011110000;
		13'd1913: color_o = 12'b000011110000;
		13'd1914: color_o = 12'b000011110000;
		13'd1915: color_o = 12'b000011110000;
		13'd1916: color_o = 12'b000011110000;
		13'd1917: color_o = 12'b000011110000;
		13'd1918: color_o = 12'b000011110000;
		13'd1919: color_o = 12'b000011110000;
		13'd1920: color_o = 12'b000011110000;
		13'd1921: color_o = 12'b000000000000;
		13'd1922: color_o = 12'b000000000000;
		13'd1923: color_o = 12'b010000000000;
		13'd1924: color_o = 12'b100000000001;
		13'd1925: color_o = 12'b100000000001;
		13'd1926: color_o = 12'b100000000001;
		13'd1927: color_o = 12'b000000000000;
		13'd1928: color_o = 12'b100000000000;
		13'd1929: color_o = 12'b100000000000;
		13'd1930: color_o = 12'b100000000000;
		13'd1931: color_o = 12'b100000000000;
		13'd1932: color_o = 12'b100000000000;
		13'd1933: color_o = 12'b000000000000;
		13'd1934: color_o = 12'b000000000000;
		13'd1935: color_o = 12'b000000000000;
		13'd1936: color_o = 12'b010000000000;
		13'd1937: color_o = 12'b010000000000;
		13'd1938: color_o = 12'b010000000000;
		13'd1939: color_o = 12'b100000000001;
		13'd1940: color_o = 12'b100000000001;
		13'd1941: color_o = 12'b100000000001;
		13'd1942: color_o = 12'b100000000000;
		13'd1943: color_o = 12'b100000000000;
		13'd1944: color_o = 12'b100000000000;
		13'd1945: color_o = 12'b100000000000;
		13'd1946: color_o = 12'b000000000000;
		13'd1947: color_o = 12'b000000000000;
		13'd1948: color_o = 12'b100000000000;
		13'd1949: color_o = 12'b100000000000;
		13'd1950: color_o = 12'b100000000000;
		13'd1951: color_o = 12'b100000000000;
		13'd1952: color_o = 12'b100000000000;
		13'd1953: color_o = 12'b100000000000;
		13'd1954: color_o = 12'b100000000000;
		13'd1955: color_o = 12'b100000000000;
		13'd1956: color_o = 12'b100000000000;
		13'd1957: color_o = 12'b000000000000;
		13'd1958: color_o = 12'b100000000001;
		13'd1959: color_o = 12'b000000000000;
		13'd1960: color_o = 12'b000000000000;
		13'd1961: color_o = 12'b011101110111;
		13'd1962: color_o = 12'b011101110111;
		13'd1963: color_o = 12'b011101110111;
		13'd1964: color_o = 12'b000000000000;
		13'd1965: color_o = 12'b100000000001;
		13'd1966: color_o = 12'b100000000001;
		13'd1967: color_o = 12'b000000000000;
		13'd1968: color_o = 12'b100000000001;
		13'd1969: color_o = 12'b000000000000;
		13'd1970: color_o = 12'b011101110111;
		13'd1971: color_o = 12'b011110011011;
		13'd1972: color_o = 12'b011110011011;
		13'd1973: color_o = 12'b011110011011;
		13'd1974: color_o = 12'b011101110111;
		13'd1975: color_o = 12'b011101110111;
		13'd1976: color_o = 12'b010001000100;
		13'd1977: color_o = 12'b000011110000;
		13'd1978: color_o = 12'b000011110000;
		13'd1979: color_o = 12'b000011110000;
		13'd1980: color_o = 12'b000011110000;
		13'd1981: color_o = 12'b000011110000;
		13'd1982: color_o = 12'b000011110000;
		13'd1983: color_o = 12'b000011110000;
		13'd1984: color_o = 12'b000011110000;
		13'd1985: color_o = 12'b000000000000;
		13'd1986: color_o = 12'b000000000000;
		13'd1987: color_o = 12'b010000000000;
		13'd1988: color_o = 12'b100000000001;
		13'd1989: color_o = 12'b100000000001;
		13'd1990: color_o = 12'b100000000001;
		13'd1991: color_o = 12'b000000000000;
		13'd1992: color_o = 12'b100000000000;
		13'd1993: color_o = 12'b000000000000;
		13'd1994: color_o = 12'b100000000000;
		13'd1995: color_o = 12'b100000000000;
		13'd1996: color_o = 12'b100000000000;
		13'd1997: color_o = 12'b100000000000;
		13'd1998: color_o = 12'b000000000000;
		13'd1999: color_o = 12'b000000000000;
		13'd2000: color_o = 12'b000000000000;
		13'd2001: color_o = 12'b000000000000;
		13'd2002: color_o = 12'b010000000000;
		13'd2003: color_o = 12'b010000000000;
		13'd2004: color_o = 12'b000000000000;
		13'd2005: color_o = 12'b000000000000;
		13'd2006: color_o = 12'b000000000000;
		13'd2007: color_o = 12'b100000000000;
		13'd2008: color_o = 12'b000000000000;
		13'd2009: color_o = 12'b000000000000;
		13'd2010: color_o = 12'b000000000000;
		13'd2011: color_o = 12'b000000000000;
		13'd2012: color_o = 12'b100000000000;
		13'd2013: color_o = 12'b100000000000;
		13'd2014: color_o = 12'b100000000000;
		13'd2015: color_o = 12'b000000000000;
		13'd2016: color_o = 12'b000000000000;
		13'd2017: color_o = 12'b000000000000;
		13'd2018: color_o = 12'b000000000000;
		13'd2019: color_o = 12'b100000000000;
		13'd2020: color_o = 12'b100000000000;
		13'd2021: color_o = 12'b000000000000;
		13'd2022: color_o = 12'b100000000001;
		13'd2023: color_o = 12'b000000000000;
		13'd2024: color_o = 12'b000000000000;
		13'd2025: color_o = 12'b011101110111;
		13'd2026: color_o = 12'b011101110111;
		13'd2027: color_o = 12'b011101110111;
		13'd2028: color_o = 12'b000000000000;
		13'd2029: color_o = 12'b100000000001;
		13'd2030: color_o = 12'b100000000001;
		13'd2031: color_o = 12'b000000000000;
		13'd2032: color_o = 12'b100000000001;
		13'd2033: color_o = 12'b100000000001;
		13'd2034: color_o = 12'b000000000000;
		13'd2035: color_o = 12'b011101110111;
		13'd2036: color_o = 12'b011101110111;
		13'd2037: color_o = 12'b011101110111;
		13'd2038: color_o = 12'b000000000000;
		13'd2039: color_o = 12'b000000000000;
		13'd2040: color_o = 12'b000000000000;
		13'd2041: color_o = 12'b000000000000;
		13'd2042: color_o = 12'b000011110000;
		13'd2043: color_o = 12'b000011110000;
		13'd2044: color_o = 12'b000011110000;
		13'd2045: color_o = 12'b000011110000;
		13'd2046: color_o = 12'b000011110000;
		13'd2047: color_o = 12'b000011110000;
		13'd2048: color_o = 12'b000011110000;
		13'd2049: color_o = 12'b000000000000;
		13'd2050: color_o = 12'b000000000000;
		13'd2051: color_o = 12'b010000000000;
		13'd2052: color_o = 12'b100000000001;
		13'd2053: color_o = 12'b100000000001;
		13'd2054: color_o = 12'b100000000001;
		13'd2055: color_o = 12'b000000000000;
		13'd2056: color_o = 12'b000000000000;
		13'd2057: color_o = 12'b000000000000;
		13'd2058: color_o = 12'b100000000001;
		13'd2059: color_o = 12'b100000000001;
		13'd2060: color_o = 12'b100000000001;
		13'd2061: color_o = 12'b100000000000;
		13'd2062: color_o = 12'b100000000000;
		13'd2063: color_o = 12'b100000000000;
		13'd2064: color_o = 12'b100000000000;
		13'd2065: color_o = 12'b000000000000;
		13'd2066: color_o = 12'b000000000000;
		13'd2067: color_o = 12'b000000000000;
		13'd2068: color_o = 12'b000000000000;
		13'd2069: color_o = 12'b100000000000;
		13'd2070: color_o = 12'b100000000001;
		13'd2071: color_o = 12'b100000000001;
		13'd2072: color_o = 12'b100000000000;
		13'd2073: color_o = 12'b000000000000;
		13'd2074: color_o = 12'b100000000000;
		13'd2075: color_o = 12'b100000000000;
		13'd2076: color_o = 12'b000000000000;
		13'd2077: color_o = 12'b000000000000;
		13'd2078: color_o = 12'b000000000000;
		13'd2079: color_o = 12'b000000000000;
		13'd2080: color_o = 12'b100000000000;
		13'd2081: color_o = 12'b100000000000;
		13'd2082: color_o = 12'b000000000000;
		13'd2083: color_o = 12'b000000000000;
		13'd2084: color_o = 12'b000000000000;
		13'd2085: color_o = 12'b000000000000;
		13'd2086: color_o = 12'b100000000001;
		13'd2087: color_o = 12'b100000000001;
		13'd2088: color_o = 12'b000000000000;
		13'd2089: color_o = 12'b000011110000;
		13'd2090: color_o = 12'b000000000000;
		13'd2091: color_o = 12'b011101110111;
		13'd2092: color_o = 12'b011101110111;
		13'd2093: color_o = 12'b011101110111;
		13'd2094: color_o = 12'b000000000000;
		13'd2095: color_o = 12'b100000000001;
		13'd2096: color_o = 12'b100000000001;
		13'd2097: color_o = 12'b000000000000;
		13'd2098: color_o = 12'b000000000000;
		13'd2099: color_o = 12'b000011110000;
		13'd2100: color_o = 12'b000011110000;
		13'd2101: color_o = 12'b000011110000;
		13'd2102: color_o = 12'b000011110000;
		13'd2103: color_o = 12'b000011110000;
		13'd2104: color_o = 12'b000011110000;
		13'd2105: color_o = 12'b000011110000;
		13'd2106: color_o = 12'b000011110000;
		13'd2107: color_o = 12'b000011110000;
		13'd2108: color_o = 12'b000011110000;
		13'd2109: color_o = 12'b000011110000;
		13'd2110: color_o = 12'b000011110000;
		13'd2111: color_o = 12'b000011110000;
		13'd2112: color_o = 12'b000011110000;
		13'd2113: color_o = 12'b000000000000;
		13'd2114: color_o = 12'b000000000000;
		13'd2115: color_o = 12'b010000000000;
		13'd2116: color_o = 12'b100000000001;
		13'd2117: color_o = 12'b100000000001;
		13'd2118: color_o = 12'b100000000001;
		13'd2119: color_o = 12'b000000000000;
		13'd2120: color_o = 12'b000000000000;
		13'd2121: color_o = 12'b100000000001;
		13'd2122: color_o = 12'b100000000001;
		13'd2123: color_o = 12'b100000000001;
		13'd2124: color_o = 12'b100000000001;
		13'd2125: color_o = 12'b100000000001;
		13'd2126: color_o = 12'b100000000000;
		13'd2127: color_o = 12'b100000000000;
		13'd2128: color_o = 12'b100000000000;
		13'd2129: color_o = 12'b100000000000;
		13'd2130: color_o = 12'b000000000000;
		13'd2131: color_o = 12'b000000000000;
		13'd2132: color_o = 12'b000000000000;
		13'd2133: color_o = 12'b010000000000;
		13'd2134: color_o = 12'b010000000000;
		13'd2135: color_o = 12'b100000000001;
		13'd2136: color_o = 12'b100000000001;
		13'd2137: color_o = 12'b100000000001;
		13'd2138: color_o = 12'b100000000000;
		13'd2139: color_o = 12'b100000000000;
		13'd2140: color_o = 12'b100000000000;
		13'd2141: color_o = 12'b100000000000;
		13'd2142: color_o = 12'b100000000000;
		13'd2143: color_o = 12'b100000000000;
		13'd2144: color_o = 12'b100000000000;
		13'd2145: color_o = 12'b000000000000;
		13'd2146: color_o = 12'b000000000000;
		13'd2147: color_o = 12'b000000000000;
		13'd2148: color_o = 12'b000000000000;
		13'd2149: color_o = 12'b000000000000;
		13'd2150: color_o = 12'b000000000000;
		13'd2151: color_o = 12'b000000000000;
		13'd2152: color_o = 12'b000011110000;
		13'd2153: color_o = 12'b000011110000;
		13'd2154: color_o = 12'b000000000000;
		13'd2155: color_o = 12'b011101110111;
		13'd2156: color_o = 12'b011101110111;
		13'd2157: color_o = 12'b011101110111;
		13'd2158: color_o = 12'b000000000000;
		13'd2159: color_o = 12'b000000000000;
		13'd2160: color_o = 12'b000000000000;
		13'd2161: color_o = 12'b000011110000;
		13'd2162: color_o = 12'b000011110000;
		13'd2163: color_o = 12'b000011110000;
		13'd2164: color_o = 12'b000011110000;
		13'd2165: color_o = 12'b000011110000;
		13'd2166: color_o = 12'b000011110000;
		13'd2167: color_o = 12'b000011110000;
		13'd2168: color_o = 12'b000011110000;
		13'd2169: color_o = 12'b000011110000;
		13'd2170: color_o = 12'b000011110000;
		13'd2171: color_o = 12'b000011110000;
		13'd2172: color_o = 12'b000011110000;
		13'd2173: color_o = 12'b000011110000;
		13'd2174: color_o = 12'b000011110000;
		13'd2175: color_o = 12'b000011110000;
		13'd2176: color_o = 12'b000011110000;
		13'd2177: color_o = 12'b000000000000;
		13'd2178: color_o = 12'b000000000000;
		13'd2179: color_o = 12'b010000000000;
		13'd2180: color_o = 12'b010000000000;
		13'd2181: color_o = 12'b100000000001;
		13'd2182: color_o = 12'b000000000000;
		13'd2183: color_o = 12'b000000000000;
		13'd2184: color_o = 12'b000000000000;
		13'd2185: color_o = 12'b000000000000;
		13'd2186: color_o = 12'b000000000000;
		13'd2187: color_o = 12'b100000000001;
		13'd2188: color_o = 12'b100000000001;
		13'd2189: color_o = 12'b100000000001;
		13'd2190: color_o = 12'b100000000001;
		13'd2191: color_o = 12'b100000000001;
		13'd2192: color_o = 12'b100000000000;
		13'd2193: color_o = 12'b100000000000;
		13'd2194: color_o = 12'b000000000000;
		13'd2195: color_o = 12'b000000000000;
		13'd2196: color_o = 12'b000000000000;
		13'd2197: color_o = 12'b000000000000;
		13'd2198: color_o = 12'b000000000000;
		13'd2199: color_o = 12'b010000000000;
		13'd2200: color_o = 12'b010000000000;
		13'd2201: color_o = 12'b010000000000;
		13'd2202: color_o = 12'b100000000001;
		13'd2203: color_o = 12'b100000000001;
		13'd2204: color_o = 12'b100000000001;
		13'd2205: color_o = 12'b100000000001;
		13'd2206: color_o = 12'b100000000001;
		13'd2207: color_o = 12'b000000000000;
		13'd2208: color_o = 12'b000000000000;
		13'd2209: color_o = 12'b000000000000;
		13'd2210: color_o = 12'b000000000000;
		13'd2211: color_o = 12'b000000000000;
		13'd2212: color_o = 12'b000000000000;
		13'd2213: color_o = 12'b000000000000;
		13'd2214: color_o = 12'b000000000000;
		13'd2215: color_o = 12'b000000000000;
		13'd2216: color_o = 12'b000011110000;
		13'd2217: color_o = 12'b000011110000;
		13'd2218: color_o = 12'b000000000000;
		13'd2219: color_o = 12'b011101110111;
		13'd2220: color_o = 12'b011101110111;
		13'd2221: color_o = 12'b000000000000;
		13'd2222: color_o = 12'b000000000000;
		13'd2223: color_o = 12'b000011110000;
		13'd2224: color_o = 12'b000011110000;
		13'd2225: color_o = 12'b000011110000;
		13'd2226: color_o = 12'b000011110000;
		13'd2227: color_o = 12'b000011110000;
		13'd2228: color_o = 12'b000011110000;
		13'd2229: color_o = 12'b000011110000;
		13'd2230: color_o = 12'b000011110000;
		13'd2231: color_o = 12'b000011110000;
		13'd2232: color_o = 12'b000011110000;
		13'd2233: color_o = 12'b000011110000;
		13'd2234: color_o = 12'b000011110000;
		13'd2235: color_o = 12'b000011110000;
		13'd2236: color_o = 12'b000011110000;
		13'd2237: color_o = 12'b000011110000;
		13'd2238: color_o = 12'b000011110000;
		13'd2239: color_o = 12'b000011110000;
		13'd2240: color_o = 12'b000011110000;
		13'd2241: color_o = 12'b000000000000;
		13'd2242: color_o = 12'b000000000000;
		13'd2243: color_o = 12'b010000000000;
		13'd2244: color_o = 12'b010000000000;
		13'd2245: color_o = 12'b000000000000;
		13'd2246: color_o = 12'b000000000000;
		13'd2247: color_o = 12'b100000000000;
		13'd2248: color_o = 12'b000000000000;
		13'd2249: color_o = 12'b000000000000;
		13'd2250: color_o = 12'b000000000000;
		13'd2251: color_o = 12'b100000000001;
		13'd2252: color_o = 12'b100000000001;
		13'd2253: color_o = 12'b100000000001;
		13'd2254: color_o = 12'b100000000001;
		13'd2255: color_o = 12'b100000000001;
		13'd2256: color_o = 12'b100000000001;
		13'd2257: color_o = 12'b100000000001;
		13'd2258: color_o = 12'b100000000000;
		13'd2259: color_o = 12'b000000000000;
		13'd2260: color_o = 12'b000000000000;
		13'd2261: color_o = 12'b000000000000;
		13'd2262: color_o = 12'b000000000000;
		13'd2263: color_o = 12'b000000000000;
		13'd2264: color_o = 12'b000000000000;
		13'd2265: color_o = 12'b000000000000;
		13'd2266: color_o = 12'b010000000000;
		13'd2267: color_o = 12'b010000000000;
		13'd2268: color_o = 12'b010000000000;
		13'd2269: color_o = 12'b010000000000;
		13'd2270: color_o = 12'b010000000000;
		13'd2271: color_o = 12'b000000000000;
		13'd2272: color_o = 12'b000011110000;
		13'd2273: color_o = 12'b000011110000;
		13'd2274: color_o = 12'b000011110000;
		13'd2275: color_o = 12'b000011110000;
		13'd2276: color_o = 12'b000011110000;
		13'd2277: color_o = 12'b000011110000;
		13'd2278: color_o = 12'b000011110000;
		13'd2279: color_o = 12'b000011110000;
		13'd2280: color_o = 12'b000011110000;
		13'd2281: color_o = 12'b000011110000;
		13'd2282: color_o = 12'b000000000000;
		13'd2283: color_o = 12'b011101110111;
		13'd2284: color_o = 12'b000000000000;
		13'd2285: color_o = 12'b000000000000;
		13'd2286: color_o = 12'b000011110000;
		13'd2287: color_o = 12'b000011110000;
		13'd2288: color_o = 12'b000011110000;
		13'd2289: color_o = 12'b000011110000;
		13'd2290: color_o = 12'b000011110000;
		13'd2291: color_o = 12'b000011110000;
		13'd2292: color_o = 12'b000011110000;
		13'd2293: color_o = 12'b000011110000;
		13'd2294: color_o = 12'b000011110000;
		13'd2295: color_o = 12'b000011110000;
		13'd2296: color_o = 12'b000011110000;
		13'd2297: color_o = 12'b000011110000;
		13'd2298: color_o = 12'b000011110000;
		13'd2299: color_o = 12'b000011110000;
		13'd2300: color_o = 12'b000011110000;
		13'd2301: color_o = 12'b000011110000;
		13'd2302: color_o = 12'b000011110000;
		13'd2303: color_o = 12'b000011110000;
		13'd2304: color_o = 12'b000011110000;
		13'd2305: color_o = 12'b000000000000;
		13'd2306: color_o = 12'b000000000000;
		13'd2307: color_o = 12'b010000000000;
		13'd2308: color_o = 12'b000000000000;
		13'd2309: color_o = 12'b000000000000;
		13'd2310: color_o = 12'b100000000000;
		13'd2311: color_o = 12'b100000000000;
		13'd2312: color_o = 12'b000000000000;
		13'd2313: color_o = 12'b000000000000;
		13'd2314: color_o = 12'b000000000000;
		13'd2315: color_o = 12'b000000000000;
		13'd2316: color_o = 12'b100000000001;
		13'd2317: color_o = 12'b100000000001;
		13'd2318: color_o = 12'b100000000001;
		13'd2319: color_o = 12'b100000000001;
		13'd2320: color_o = 12'b100000000000;
		13'd2321: color_o = 12'b100000000001;
		13'd2322: color_o = 12'b100000000001;
		13'd2323: color_o = 12'b100000000001;
		13'd2324: color_o = 12'b100000000000;
		13'd2325: color_o = 12'b100000000000;
		13'd2326: color_o = 12'b100000000000;
		13'd2327: color_o = 12'b000000000000;
		13'd2328: color_o = 12'b000000000000;
		13'd2329: color_o = 12'b000000000000;
		13'd2330: color_o = 12'b000000000000;
		13'd2331: color_o = 12'b000000000000;
		13'd2332: color_o = 12'b000000000000;
		13'd2333: color_o = 12'b000000000000;
		13'd2334: color_o = 12'b000000000000;
		13'd2335: color_o = 12'b000011110000;
		13'd2336: color_o = 12'b000011110000;
		13'd2337: color_o = 12'b000011110000;
		13'd2338: color_o = 12'b000011110000;
		13'd2339: color_o = 12'b000011110000;
		13'd2340: color_o = 12'b000011110000;
		13'd2341: color_o = 12'b000011110000;
		13'd2342: color_o = 12'b000011110000;
		13'd2343: color_o = 12'b000011110000;
		13'd2344: color_o = 12'b000011110000;
		13'd2345: color_o = 12'b000011110000;
		13'd2346: color_o = 12'b000000000000;
		13'd2347: color_o = 12'b000000000000;
		13'd2348: color_o = 12'b000011110000;
		13'd2349: color_o = 12'b000011110000;
		13'd2350: color_o = 12'b000011110000;
		13'd2351: color_o = 12'b000011110000;
		13'd2352: color_o = 12'b000011110000;
		13'd2353: color_o = 12'b000011110000;
		13'd2354: color_o = 12'b000011110000;
		13'd2355: color_o = 12'b000011110000;
		13'd2356: color_o = 12'b000011110000;
		13'd2357: color_o = 12'b000011110000;
		13'd2358: color_o = 12'b000011110000;
		13'd2359: color_o = 12'b000011110000;
		13'd2360: color_o = 12'b000011110000;
		13'd2361: color_o = 12'b000011110000;
		13'd2362: color_o = 12'b000011110000;
		13'd2363: color_o = 12'b000011110000;
		13'd2364: color_o = 12'b000011110000;
		13'd2365: color_o = 12'b000011110000;
		13'd2366: color_o = 12'b000011110000;
		13'd2367: color_o = 12'b000011110000;
		13'd2368: color_o = 12'b000011110000;
		13'd2369: color_o = 12'b000000000000;
		13'd2370: color_o = 12'b000000000000;
		13'd2371: color_o = 12'b000000000000;
		13'd2372: color_o = 12'b000000000000;
		13'd2373: color_o = 12'b000000000000;
		13'd2374: color_o = 12'b100000000001;
		13'd2375: color_o = 12'b100000000001;
		13'd2376: color_o = 12'b000000000000;
		13'd2377: color_o = 12'b000000000000;
		13'd2378: color_o = 12'b100000000000;
		13'd2379: color_o = 12'b000000000000;
		13'd2380: color_o = 12'b000000000000;
		13'd2381: color_o = 12'b000000000000;
		13'd2382: color_o = 12'b000000000000;
		13'd2383: color_o = 12'b100000000000;
		13'd2384: color_o = 12'b100000000001;
		13'd2385: color_o = 12'b100000000001;
		13'd2386: color_o = 12'b100000000001;
		13'd2387: color_o = 12'b100000000001;
		13'd2388: color_o = 12'b100000000001;
		13'd2389: color_o = 12'b100000000000;
		13'd2390: color_o = 12'b100000000000;
		13'd2391: color_o = 12'b100000000000;
		13'd2392: color_o = 12'b000000000000;
		13'd2393: color_o = 12'b000000000000;
		13'd2394: color_o = 12'b100000000000;
		13'd2395: color_o = 12'b100000000000;
		13'd2396: color_o = 12'b100000000000;
		13'd2397: color_o = 12'b000000000000;
		13'd2398: color_o = 12'b000000000000;
		13'd2399: color_o = 12'b000011110000;
		13'd2400: color_o = 12'b000011110000;
		13'd2401: color_o = 12'b000011110000;
		13'd2402: color_o = 12'b000011110000;
		13'd2403: color_o = 12'b000011110000;
		13'd2404: color_o = 12'b000011110000;
		13'd2405: color_o = 12'b000011110000;
		13'd2406: color_o = 12'b000011110000;
		13'd2407: color_o = 12'b000011110000;
		13'd2408: color_o = 12'b000011110000;
		13'd2409: color_o = 12'b000011110000;
		13'd2410: color_o = 12'b000000000000;
		13'd2411: color_o = 12'b000011110000;
		13'd2412: color_o = 12'b000011110000;
		13'd2413: color_o = 12'b000011110000;
		13'd2414: color_o = 12'b000011110000;
		13'd2415: color_o = 12'b000011110000;
		13'd2416: color_o = 12'b000011110000;
		13'd2417: color_o = 12'b000011110000;
		13'd2418: color_o = 12'b000011110000;
		13'd2419: color_o = 12'b000011110000;
		13'd2420: color_o = 12'b000011110000;
		13'd2421: color_o = 12'b000011110000;
		13'd2422: color_o = 12'b000011110000;
		13'd2423: color_o = 12'b000011110000;
		13'd2424: color_o = 12'b000011110000;
		13'd2425: color_o = 12'b000011110000;
		13'd2426: color_o = 12'b000011110000;
		13'd2427: color_o = 12'b000011110000;
		13'd2428: color_o = 12'b000011110000;
		13'd2429: color_o = 12'b000011110000;
		13'd2430: color_o = 12'b000011110000;
		13'd2431: color_o = 12'b000011110000;
		13'd2432: color_o = 12'b000011110000;
		13'd2433: color_o = 12'b000011110000;
		13'd2434: color_o = 12'b000011110000;
		13'd2435: color_o = 12'b000011110000;
		13'd2436: color_o = 12'b000000000000;
		13'd2437: color_o = 12'b000000000000;
		13'd2438: color_o = 12'b000000000000;
		13'd2439: color_o = 12'b000000000000;
		13'd2440: color_o = 12'b000000000000;
		13'd2441: color_o = 12'b000000000000;
		13'd2442: color_o = 12'b000000000000;
		13'd2443: color_o = 12'b000000000000;
		13'd2444: color_o = 12'b100000000000;
		13'd2445: color_o = 12'b000000000000;
		13'd2446: color_o = 12'b000000000000;
		13'd2447: color_o = 12'b000000000000;
		13'd2448: color_o = 12'b000000000000;
		13'd2449: color_o = 12'b000000000000;
		13'd2450: color_o = 12'b000000000000;
		13'd2451: color_o = 12'b000000000000;
		13'd2452: color_o = 12'b100000000001;
		13'd2453: color_o = 12'b100000000001;
		13'd2454: color_o = 12'b000000000000;
		13'd2455: color_o = 12'b000000000000;
		13'd2456: color_o = 12'b000000000000;
		13'd2457: color_o = 12'b000000000000;
		13'd2458: color_o = 12'b000000000000;
		13'd2459: color_o = 12'b000000000000;
		13'd2460: color_o = 12'b000000000000;
		13'd2461: color_o = 12'b000000000000;
		13'd2462: color_o = 12'b000011110000;
		13'd2463: color_o = 12'b000011110000;
		13'd2464: color_o = 12'b000011110000;
		13'd2465: color_o = 12'b000011110000;
		13'd2466: color_o = 12'b000011110000;
		13'd2467: color_o = 12'b000011110000;
		13'd2468: color_o = 12'b000011110000;
		13'd2469: color_o = 12'b000011110000;
		13'd2470: color_o = 12'b000011110000;
		13'd2471: color_o = 12'b000011110000;
		13'd2472: color_o = 12'b000011110000;
		13'd2473: color_o = 12'b000011110000;
		13'd2474: color_o = 12'b000011110000;
		13'd2475: color_o = 12'b000011110000;
		13'd2476: color_o = 12'b000011110000;
		13'd2477: color_o = 12'b000011110000;
		13'd2478: color_o = 12'b000011110000;
		13'd2479: color_o = 12'b000011110000;
		13'd2480: color_o = 12'b000011110000;
		13'd2481: color_o = 12'b000011110000;
		13'd2482: color_o = 12'b000011110000;
		13'd2483: color_o = 12'b000011110000;
		13'd2484: color_o = 12'b000011110000;
		13'd2485: color_o = 12'b000011110000;
		13'd2486: color_o = 12'b000011110000;
		13'd2487: color_o = 12'b000011110000;
		13'd2488: color_o = 12'b000011110000;
		13'd2489: color_o = 12'b000011110000;
		13'd2490: color_o = 12'b000011110000;
		13'd2491: color_o = 12'b000011110000;
		13'd2492: color_o = 12'b000011110000;
		13'd2493: color_o = 12'b000011110000;
		13'd2494: color_o = 12'b000011110000;
		13'd2495: color_o = 12'b000011110000;
		13'd2496: color_o = 12'b000011110000;
		13'd2497: color_o = 12'b000011110000;
		13'd2498: color_o = 12'b000011110000;
		13'd2499: color_o = 12'b000011110000;
		13'd2500: color_o = 12'b000011110000;
		13'd2501: color_o = 12'b000011110000;
		13'd2502: color_o = 12'b000000000000;
		13'd2503: color_o = 12'b000000000000;
		13'd2504: color_o = 12'b000000000000;
		13'd2505: color_o = 12'b000000000000;
		13'd2506: color_o = 12'b000000000000;
		13'd2507: color_o = 12'b000000000000;
		13'd2508: color_o = 12'b100000000000;
		13'd2509: color_o = 12'b100000000000;
		13'd2510: color_o = 12'b100000000000;
		13'd2511: color_o = 12'b100000000000;
		13'd2512: color_o = 12'b100000000000;
		13'd2513: color_o = 12'b100000000000;
		13'd2514: color_o = 12'b100000000000;
		13'd2515: color_o = 12'b000000000000;
		13'd2516: color_o = 12'b000000000000;
		13'd2517: color_o = 12'b000000000000;
		13'd2518: color_o = 12'b000000000000;
		13'd2519: color_o = 12'b000000000000;
		13'd2520: color_o = 12'b000000000000;
		13'd2521: color_o = 12'b000000000000;
		13'd2522: color_o = 12'b000000000000;
		13'd2523: color_o = 12'b000000000000;
		13'd2524: color_o = 12'b000000000000;
		13'd2525: color_o = 12'b000011110000;
		13'd2526: color_o = 12'b000011110000;
		13'd2527: color_o = 12'b000011110000;
		13'd2528: color_o = 12'b000011110000;
		13'd2529: color_o = 12'b000011110000;
		13'd2530: color_o = 12'b000011110000;
		13'd2531: color_o = 12'b000011110000;
		13'd2532: color_o = 12'b000011110000;
		13'd2533: color_o = 12'b000011110000;
		13'd2534: color_o = 12'b000011110000;
		13'd2535: color_o = 12'b000011110000;
		13'd2536: color_o = 12'b000011110000;
		13'd2537: color_o = 12'b000011110000;
		13'd2538: color_o = 12'b000011110000;
		13'd2539: color_o = 12'b000011110000;
		13'd2540: color_o = 12'b000011110000;
		13'd2541: color_o = 12'b000011110000;
		13'd2542: color_o = 12'b000011110000;
		13'd2543: color_o = 12'b000011110000;
		13'd2544: color_o = 12'b000011110000;
		13'd2545: color_o = 12'b000011110000;
		13'd2546: color_o = 12'b000011110000;
		13'd2547: color_o = 12'b000011110000;
		13'd2548: color_o = 12'b000011110000;
		13'd2549: color_o = 12'b000011110000;
		13'd2550: color_o = 12'b000011110000;
		13'd2551: color_o = 12'b000011110000;
		13'd2552: color_o = 12'b000011110000;
		13'd2553: color_o = 12'b000011110000;
		13'd2554: color_o = 12'b000011110000;
		13'd2555: color_o = 12'b000011110000;
		13'd2556: color_o = 12'b000011110000;
		13'd2557: color_o = 12'b000011110000;
		13'd2558: color_o = 12'b000011110000;
		13'd2559: color_o = 12'b000011110000;
		13'd2560: color_o = 12'b000011110000;
		13'd2561: color_o = 12'b000011110000;
		13'd2562: color_o = 12'b000011110000;
		13'd2563: color_o = 12'b000011110000;
		13'd2564: color_o = 12'b000011110000;
		13'd2565: color_o = 12'b000011110000;
		13'd2566: color_o = 12'b000011110000;
		13'd2567: color_o = 12'b000011110000;
		13'd2568: color_o = 12'b000011110000;
		13'd2569: color_o = 12'b000011110000;
		13'd2570: color_o = 12'b000011110000;
		13'd2571: color_o = 12'b000011110000;
		13'd2572: color_o = 12'b000011110000;
		13'd2573: color_o = 12'b000011110000;
		13'd2574: color_o = 12'b000011110000;
		13'd2575: color_o = 12'b000011110000;
		13'd2576: color_o = 12'b000011110000;
		13'd2577: color_o = 12'b000011110000;
		13'd2578: color_o = 12'b000011110000;
		13'd2579: color_o = 12'b000011110000;
		13'd2580: color_o = 12'b000011110000;
		13'd2581: color_o = 12'b000011110000;
		13'd2582: color_o = 12'b000011110000;
		13'd2583: color_o = 12'b000011110000;
		13'd2584: color_o = 12'b000011110000;
		13'd2585: color_o = 12'b000011110000;
		13'd2586: color_o = 12'b000011110000;
		13'd2587: color_o = 12'b000011110000;
		13'd2588: color_o = 12'b000011110000;
		13'd2589: color_o = 12'b000011110000;
		13'd2590: color_o = 12'b000011110000;
		13'd2591: color_o = 12'b000011110000;
		13'd2592: color_o = 12'b000011110000;
		13'd2593: color_o = 12'b000011110000;
		13'd2594: color_o = 12'b000011110000;
		13'd2595: color_o = 12'b000011110000;
		13'd2596: color_o = 12'b000011110000;
		13'd2597: color_o = 12'b000011110000;
		13'd2598: color_o = 12'b000011110000;
		13'd2599: color_o = 12'b000011110000;
		13'd2600: color_o = 12'b000011110000;
		13'd2601: color_o = 12'b000011110000;
		13'd2602: color_o = 12'b000011110000;
		13'd2603: color_o = 12'b000011110000;
		13'd2604: color_o = 12'b000011110000;
		13'd2605: color_o = 12'b000011110000;
		13'd2606: color_o = 12'b000011110000;
		13'd2607: color_o = 12'b000011110000;
		13'd2608: color_o = 12'b000011110000;
		13'd2609: color_o = 12'b000011110000;
		13'd2610: color_o = 12'b000011110000;
		13'd2611: color_o = 12'b000011110000;
		13'd2612: color_o = 12'b000011110000;
		13'd2613: color_o = 12'b000011110000;
		13'd2614: color_o = 12'b000011110000;
		13'd2615: color_o = 12'b000011110000;
		13'd2616: color_o = 12'b000011110000;
		13'd2617: color_o = 12'b000011110000;
		13'd2618: color_o = 12'b000011110000;
		13'd2619: color_o = 12'b000011110000;
		13'd2620: color_o = 12'b000011110000;
		13'd2621: color_o = 12'b000011110000;
		13'd2622: color_o = 12'b000011110000;
		13'd2623: color_o = 12'b000011110000;
		13'd2624: color_o = 12'b000011110000;
		13'd2625: color_o = 12'b000011110000;
		13'd2626: color_o = 12'b000011110000;
		13'd2627: color_o = 12'b000011110000;
		13'd2628: color_o = 12'b000011110000;
		13'd2629: color_o = 12'b000011110000;
		13'd2630: color_o = 12'b000011110000;
		13'd2631: color_o = 12'b000011110000;
		13'd2632: color_o = 12'b000011110000;
		13'd2633: color_o = 12'b000011110000;
		13'd2634: color_o = 12'b000011110000;
		13'd2635: color_o = 12'b000011110000;
		13'd2636: color_o = 12'b000011110000;
		13'd2637: color_o = 12'b000011110000;
		13'd2638: color_o = 12'b000011110000;
		13'd2639: color_o = 12'b000011110000;
		13'd2640: color_o = 12'b000011110000;
		13'd2641: color_o = 12'b000011110000;
		13'd2642: color_o = 12'b000011110000;
		13'd2643: color_o = 12'b000011110000;
		13'd2644: color_o = 12'b000011110000;
		13'd2645: color_o = 12'b000011110000;
		13'd2646: color_o = 12'b000011110000;
		13'd2647: color_o = 12'b000011110000;
		13'd2648: color_o = 12'b000011110000;
		13'd2649: color_o = 12'b000011110000;
		13'd2650: color_o = 12'b000011110000;
		13'd2651: color_o = 12'b000011110000;
		13'd2652: color_o = 12'b000011110000;
		13'd2653: color_o = 12'b000011110000;
		13'd2654: color_o = 12'b000011110000;
		13'd2655: color_o = 12'b000011110000;
		13'd2656: color_o = 12'b000011110000;
		13'd2657: color_o = 12'b000011110000;
		13'd2658: color_o = 12'b000011110000;
		13'd2659: color_o = 12'b000011110000;
		13'd2660: color_o = 12'b000011110000;
		13'd2661: color_o = 12'b000011110000;
		13'd2662: color_o = 12'b000011110000;
		13'd2663: color_o = 12'b000011110000;
		13'd2664: color_o = 12'b000011110000;
		13'd2665: color_o = 12'b000011110000;
		13'd2666: color_o = 12'b000011110000;
		13'd2667: color_o = 12'b000011110000;
		13'd2668: color_o = 12'b000011110000;
		13'd2669: color_o = 12'b000011110000;
		13'd2670: color_o = 12'b000011110000;
		13'd2671: color_o = 12'b000011110000;
		13'd2672: color_o = 12'b000011110000;
		13'd2673: color_o = 12'b000011110000;
		13'd2674: color_o = 12'b000011110000;
		13'd2675: color_o = 12'b000011110000;
		13'd2676: color_o = 12'b000011110000;
		13'd2677: color_o = 12'b000011110000;
		13'd2678: color_o = 12'b000011110000;
		13'd2679: color_o = 12'b000011110000;
		13'd2680: color_o = 12'b000011110000;
		13'd2681: color_o = 12'b000011110000;
		13'd2682: color_o = 12'b000011110000;
		13'd2683: color_o = 12'b000011110000;
		13'd2684: color_o = 12'b000011110000;
		13'd2685: color_o = 12'b000011110000;
		13'd2686: color_o = 12'b000011110000;
		13'd2687: color_o = 12'b000011110000;
		13'd2688: color_o = 12'b000011110000;
		13'd2689: color_o = 12'b000011110000;
		13'd2690: color_o = 12'b000011110000;
		13'd2691: color_o = 12'b000011110000;
		13'd2692: color_o = 12'b000011110000;
		13'd2693: color_o = 12'b000011110000;
		13'd2694: color_o = 12'b000011110000;
		13'd2695: color_o = 12'b000011110000;
		13'd2696: color_o = 12'b000011110000;
		13'd2697: color_o = 12'b000011110000;
		13'd2698: color_o = 12'b000011110000;
		13'd2699: color_o = 12'b000011110000;
		13'd2700: color_o = 12'b000011110000;
		13'd2701: color_o = 12'b000011110000;
		13'd2702: color_o = 12'b000011110000;
		13'd2703: color_o = 12'b000011110000;
		13'd2704: color_o = 12'b000011110000;
		13'd2705: color_o = 12'b000011110000;
		13'd2706: color_o = 12'b000011110000;
		13'd2707: color_o = 12'b000011110000;
		13'd2708: color_o = 12'b000011110000;
		13'd2709: color_o = 12'b000011110000;
		13'd2710: color_o = 12'b000011110000;
		13'd2711: color_o = 12'b000011110000;
		13'd2712: color_o = 12'b000011110000;
		13'd2713: color_o = 12'b000011110000;
		13'd2714: color_o = 12'b000011110000;
		13'd2715: color_o = 12'b000011110000;
		13'd2716: color_o = 12'b000011110000;
		13'd2717: color_o = 12'b000011110000;
		13'd2718: color_o = 12'b000011110000;
		13'd2719: color_o = 12'b000011110000;
		13'd2720: color_o = 12'b000011110000;
		13'd2721: color_o = 12'b000011110000;
		13'd2722: color_o = 12'b000011110000;
		13'd2723: color_o = 12'b000011110000;
		13'd2724: color_o = 12'b000011110000;
		13'd2725: color_o = 12'b000011110000;
		13'd2726: color_o = 12'b000011110000;
		13'd2727: color_o = 12'b000011110000;
		13'd2728: color_o = 12'b000011110000;
		13'd2729: color_o = 12'b000011110000;
		13'd2730: color_o = 12'b000011110000;
		13'd2731: color_o = 12'b000011110000;
		13'd2732: color_o = 12'b000011110000;
		13'd2733: color_o = 12'b000011110000;
		13'd2734: color_o = 12'b000011110000;
		13'd2735: color_o = 12'b000011110000;
		13'd2736: color_o = 12'b000011110000;
		13'd2737: color_o = 12'b000011110000;
		13'd2738: color_o = 12'b000011110000;
		13'd2739: color_o = 12'b000011110000;
		13'd2740: color_o = 12'b000011110000;
		13'd2741: color_o = 12'b000011110000;
		13'd2742: color_o = 12'b000011110000;
		13'd2743: color_o = 12'b000011110000;
		13'd2744: color_o = 12'b000011110000;
		13'd2745: color_o = 12'b000011110000;
		13'd2746: color_o = 12'b000011110000;
		13'd2747: color_o = 12'b000011110000;
		13'd2748: color_o = 12'b000011110000;
		13'd2749: color_o = 12'b000011110000;
		13'd2750: color_o = 12'b000011110000;
		13'd2751: color_o = 12'b000011110000;
		13'd2752: color_o = 12'b000011110000;
		13'd2753: color_o = 12'b000011110000;
		13'd2754: color_o = 12'b000011110000;
		13'd2755: color_o = 12'b000011110000;
		13'd2756: color_o = 12'b000011110000;
		13'd2757: color_o = 12'b000011110000;
		13'd2758: color_o = 12'b000011110000;
		13'd2759: color_o = 12'b000011110000;
		13'd2760: color_o = 12'b000011110000;
		13'd2761: color_o = 12'b000011110000;
		13'd2762: color_o = 12'b000011110000;
		13'd2763: color_o = 12'b000011110000;
		13'd2764: color_o = 12'b000011110000;
		13'd2765: color_o = 12'b000011110000;
		13'd2766: color_o = 12'b000011110000;
		13'd2767: color_o = 12'b000011110000;
		13'd2768: color_o = 12'b000011110000;
		13'd2769: color_o = 12'b000011110000;
		13'd2770: color_o = 12'b000011110000;
		13'd2771: color_o = 12'b000011110000;
		13'd2772: color_o = 12'b000011110000;
		13'd2773: color_o = 12'b000011110000;
		13'd2774: color_o = 12'b000011110000;
		13'd2775: color_o = 12'b000011110000;
		13'd2776: color_o = 12'b000011110000;
		13'd2777: color_o = 12'b000011110000;
		13'd2778: color_o = 12'b000011110000;
		13'd2779: color_o = 12'b000011110000;
		13'd2780: color_o = 12'b000011110000;
		13'd2781: color_o = 12'b000011110000;
		13'd2782: color_o = 12'b000011110000;
		13'd2783: color_o = 12'b000011110000;
		13'd2784: color_o = 12'b000011110000;
		13'd2785: color_o = 12'b000011110000;
		13'd2786: color_o = 12'b000011110000;
		13'd2787: color_o = 12'b000011110000;
		13'd2788: color_o = 12'b000011110000;
		13'd2789: color_o = 12'b000011110000;
		13'd2790: color_o = 12'b000011110000;
		13'd2791: color_o = 12'b000011110000;
		13'd2792: color_o = 12'b000011110000;
		13'd2793: color_o = 12'b000011110000;
		13'd2794: color_o = 12'b000011110000;
		13'd2795: color_o = 12'b000011110000;
		13'd2796: color_o = 12'b000011110000;
		13'd2797: color_o = 12'b000011110000;
		13'd2798: color_o = 12'b000011110000;
		13'd2799: color_o = 12'b000011110000;
		13'd2800: color_o = 12'b000011110000;
		13'd2801: color_o = 12'b000011110000;
		13'd2802: color_o = 12'b000011110000;
		13'd2803: color_o = 12'b000011110000;
		13'd2804: color_o = 12'b000011110000;
		13'd2805: color_o = 12'b000011110000;
		13'd2806: color_o = 12'b000011110000;
		13'd2807: color_o = 12'b000011110000;
		13'd2808: color_o = 12'b000011110000;
		13'd2809: color_o = 12'b000011110000;
		13'd2810: color_o = 12'b000011110000;
		13'd2811: color_o = 12'b000011110000;
		13'd2812: color_o = 12'b000011110000;
		13'd2813: color_o = 12'b000011110000;
		13'd2814: color_o = 12'b000011110000;
		13'd2815: color_o = 12'b000011110000;
		13'd2816: color_o = 12'b000011110000;
		13'd2817: color_o = 12'b000011110000;
		13'd2818: color_o = 12'b000011110000;
		13'd2819: color_o = 12'b000011110000;
		13'd2820: color_o = 12'b000011110000;
		13'd2821: color_o = 12'b000011110000;
		13'd2822: color_o = 12'b000011110000;
		13'd2823: color_o = 12'b000011110000;
		13'd2824: color_o = 12'b000011110000;
		13'd2825: color_o = 12'b000011110000;
		13'd2826: color_o = 12'b000011110000;
		13'd2827: color_o = 12'b000011110000;
		13'd2828: color_o = 12'b000011110000;
		13'd2829: color_o = 12'b000011110000;
		13'd2830: color_o = 12'b000011110000;
		13'd2831: color_o = 12'b000011110000;
		13'd2832: color_o = 12'b000011110000;
		13'd2833: color_o = 12'b000011110000;
		13'd2834: color_o = 12'b000011110000;
		13'd2835: color_o = 12'b000011110000;
		13'd2836: color_o = 12'b000011110000;
		13'd2837: color_o = 12'b000011110000;
		13'd2838: color_o = 12'b000011110000;
		13'd2839: color_o = 12'b000011110000;
		13'd2840: color_o = 12'b000011110000;
		13'd2841: color_o = 12'b000011110000;
		13'd2842: color_o = 12'b000011110000;
		13'd2843: color_o = 12'b000011110000;
		13'd2844: color_o = 12'b000011110000;
		13'd2845: color_o = 12'b000011110000;
		13'd2846: color_o = 12'b000011110000;
		13'd2847: color_o = 12'b000011110000;
		13'd2848: color_o = 12'b000011110000;
		13'd2849: color_o = 12'b000011110000;
		13'd2850: color_o = 12'b000011110000;
		13'd2851: color_o = 12'b000011110000;
		13'd2852: color_o = 12'b000011110000;
		13'd2853: color_o = 12'b000011110000;
		13'd2854: color_o = 12'b000011110000;
		13'd2855: color_o = 12'b000011110000;
		13'd2856: color_o = 12'b000011110000;
		13'd2857: color_o = 12'b000011110000;
		13'd2858: color_o = 12'b000011110000;
		13'd2859: color_o = 12'b000011110000;
		13'd2860: color_o = 12'b000011110000;
		13'd2861: color_o = 12'b000011110000;
		13'd2862: color_o = 12'b000011110000;
		13'd2863: color_o = 12'b000011110000;
		13'd2864: color_o = 12'b000011110000;
		13'd2865: color_o = 12'b000011110000;
		13'd2866: color_o = 12'b000011110000;
		13'd2867: color_o = 12'b000011110000;
		13'd2868: color_o = 12'b000011110000;
		13'd2869: color_o = 12'b000011110000;
		13'd2870: color_o = 12'b000011110000;
		13'd2871: color_o = 12'b000011110000;
		13'd2872: color_o = 12'b000011110000;
		13'd2873: color_o = 12'b000011110000;
		13'd2874: color_o = 12'b000011110000;
		13'd2875: color_o = 12'b000011110000;
		13'd2876: color_o = 12'b000011110000;
		13'd2877: color_o = 12'b000011110000;
		13'd2878: color_o = 12'b000011110000;
		13'd2879: color_o = 12'b000011110000;
		13'd2880: color_o = 12'b000011110000;
		13'd2881: color_o = 12'b000011110000;
		13'd2882: color_o = 12'b000011110000;
		13'd2883: color_o = 12'b000011110000;
		13'd2884: color_o = 12'b000011110000;
		13'd2885: color_o = 12'b000011110000;
		13'd2886: color_o = 12'b000011110000;
		13'd2887: color_o = 12'b000011110000;
		13'd2888: color_o = 12'b000011110000;
		13'd2889: color_o = 12'b000011110000;
		13'd2890: color_o = 12'b000011110000;
		13'd2891: color_o = 12'b000011110000;
		13'd2892: color_o = 12'b000011110000;
		13'd2893: color_o = 12'b000011110000;
		13'd2894: color_o = 12'b000000000000;
		13'd2895: color_o = 12'b000000000000;
		13'd2896: color_o = 12'b000000000000;
		13'd2897: color_o = 12'b011000000000;
		13'd2898: color_o = 12'b011000000000;
		13'd2899: color_o = 12'b011000000000;
		13'd2900: color_o = 12'b000011110000;
		13'd2901: color_o = 12'b000011110000;
		13'd2902: color_o = 12'b000011110000;
		13'd2903: color_o = 12'b000011110000;
		13'd2904: color_o = 12'b000011110000;
		13'd2905: color_o = 12'b000011110000;
		13'd2906: color_o = 12'b000011110000;
		13'd2907: color_o = 12'b000011110000;
		13'd2908: color_o = 12'b000011110000;
		13'd2909: color_o = 12'b000011110000;
		13'd2910: color_o = 12'b000011110000;
		13'd2911: color_o = 12'b000011110000;
		13'd2912: color_o = 12'b000011110000;
		13'd2913: color_o = 12'b000011110000;
		13'd2914: color_o = 12'b000011110000;
		13'd2915: color_o = 12'b000011110000;
		13'd2916: color_o = 12'b000011110000;
		13'd2917: color_o = 12'b000011110000;
		13'd2918: color_o = 12'b000011110000;
		13'd2919: color_o = 12'b000011110000;
		13'd2920: color_o = 12'b000011110000;
		13'd2921: color_o = 12'b000011110000;
		13'd2922: color_o = 12'b000011110000;
		13'd2923: color_o = 12'b000011110000;
		13'd2924: color_o = 12'b000011110000;
		13'd2925: color_o = 12'b000011110000;
		13'd2926: color_o = 12'b000011110000;
		13'd2927: color_o = 12'b000011110000;
		13'd2928: color_o = 12'b000011110000;
		13'd2929: color_o = 12'b000011110000;
		13'd2930: color_o = 12'b000011110000;
		13'd2931: color_o = 12'b000011110000;
		13'd2932: color_o = 12'b000011110000;
		13'd2933: color_o = 12'b000011110000;
		13'd2934: color_o = 12'b000011110000;
		13'd2935: color_o = 12'b000011110000;
		13'd2936: color_o = 12'b000011110000;
		13'd2937: color_o = 12'b000011110000;
		13'd2938: color_o = 12'b000011110000;
		13'd2939: color_o = 12'b000011110000;
		13'd2940: color_o = 12'b000011110000;
		13'd2941: color_o = 12'b000011110000;
		13'd2942: color_o = 12'b000011110000;
		13'd2943: color_o = 12'b000011110000;
		13'd2944: color_o = 12'b000011110000;
		13'd2945: color_o = 12'b000011110000;
		13'd2946: color_o = 12'b000011110000;
		13'd2947: color_o = 12'b000011110000;
		13'd2948: color_o = 12'b000011110000;
		13'd2949: color_o = 12'b000011110000;
		13'd2950: color_o = 12'b000011110000;
		13'd2951: color_o = 12'b000011110000;
		13'd2952: color_o = 12'b000011110000;
		13'd2953: color_o = 12'b000011110000;
		13'd2954: color_o = 12'b000011110000;
		13'd2955: color_o = 12'b000011110000;
		13'd2956: color_o = 12'b000011110000;
		13'd2957: color_o = 12'b000000000000;
		13'd2958: color_o = 12'b000000000000;
		13'd2959: color_o = 12'b000000000000;
		13'd2960: color_o = 12'b100000000000;
		13'd2961: color_o = 12'b011000000000;
		13'd2962: color_o = 12'b011000000000;
		13'd2963: color_o = 12'b011000000000;
		13'd2964: color_o = 12'b011000000000;
		13'd2965: color_o = 12'b011000000000;
		13'd2966: color_o = 12'b011000000000;
		13'd2967: color_o = 12'b011000000000;
		13'd2968: color_o = 12'b000011110000;
		13'd2969: color_o = 12'b000011110000;
		13'd2970: color_o = 12'b000011110000;
		13'd2971: color_o = 12'b000011110000;
		13'd2972: color_o = 12'b000011110000;
		13'd2973: color_o = 12'b000011110000;
		13'd2974: color_o = 12'b000011110000;
		13'd2975: color_o = 12'b000011110000;
		13'd2976: color_o = 12'b000011110000;
		13'd2977: color_o = 12'b000011110000;
		13'd2978: color_o = 12'b000011110000;
		13'd2979: color_o = 12'b000011110000;
		13'd2980: color_o = 12'b000011110000;
		13'd2981: color_o = 12'b000011110000;
		13'd2982: color_o = 12'b000011110000;
		13'd2983: color_o = 12'b000011110000;
		13'd2984: color_o = 12'b000011110000;
		13'd2985: color_o = 12'b000011110000;
		13'd2986: color_o = 12'b000011110000;
		13'd2987: color_o = 12'b000011110000;
		13'd2988: color_o = 12'b000011110000;
		13'd2989: color_o = 12'b000011110000;
		13'd2990: color_o = 12'b000011110000;
		13'd2991: color_o = 12'b000011110000;
		13'd2992: color_o = 12'b000011110000;
		13'd2993: color_o = 12'b000011110000;
		13'd2994: color_o = 12'b000011110000;
		13'd2995: color_o = 12'b000011110000;
		13'd2996: color_o = 12'b000011110000;
		13'd2997: color_o = 12'b000011110000;
		13'd2998: color_o = 12'b000011110000;
		13'd2999: color_o = 12'b000011110000;
		13'd3000: color_o = 12'b000011110000;
		13'd3001: color_o = 12'b000011110000;
		13'd3002: color_o = 12'b000011110000;
		13'd3003: color_o = 12'b000011110000;
		13'd3004: color_o = 12'b000011110000;
		13'd3005: color_o = 12'b000011110000;
		13'd3006: color_o = 12'b000011110000;
		13'd3007: color_o = 12'b000011110000;
		13'd3008: color_o = 12'b000011110000;
		13'd3009: color_o = 12'b000011110000;
		13'd3010: color_o = 12'b000011110000;
		13'd3011: color_o = 12'b000011110000;
		13'd3012: color_o = 12'b000011110000;
		13'd3013: color_o = 12'b000011110000;
		13'd3014: color_o = 12'b000011110000;
		13'd3015: color_o = 12'b000011110000;
		13'd3016: color_o = 12'b000011110000;
		13'd3017: color_o = 12'b000011110000;
		13'd3018: color_o = 12'b000011110000;
		13'd3019: color_o = 12'b000000000000;
		13'd3020: color_o = 12'b000000000000;
		13'd3021: color_o = 12'b000000000000;
		13'd3022: color_o = 12'b100000000000;
		13'd3023: color_o = 12'b100000000000;
		13'd3024: color_o = 12'b100000000000;
		13'd3025: color_o = 12'b100000000000;
		13'd3026: color_o = 12'b100000000000;
		13'd3027: color_o = 12'b100000000000;
		13'd3028: color_o = 12'b011000000000;
		13'd3029: color_o = 12'b011000000000;
		13'd3030: color_o = 12'b100000000000;
		13'd3031: color_o = 12'b011000000000;
		13'd3032: color_o = 12'b011000000000;
		13'd3033: color_o = 12'b011000000000;
		13'd3034: color_o = 12'b011000000000;
		13'd3035: color_o = 12'b011000000000;
		13'd3036: color_o = 12'b011000000000;
		13'd3037: color_o = 12'b000011110000;
		13'd3038: color_o = 12'b000011110000;
		13'd3039: color_o = 12'b000011110000;
		13'd3040: color_o = 12'b000011110000;
		13'd3041: color_o = 12'b000011110000;
		13'd3042: color_o = 12'b000011110000;
		13'd3043: color_o = 12'b000011110000;
		13'd3044: color_o = 12'b000011110000;
		13'd3045: color_o = 12'b000011110000;
		13'd3046: color_o = 12'b000011110000;
		13'd3047: color_o = 12'b000011110000;
		13'd3048: color_o = 12'b000011110000;
		13'd3049: color_o = 12'b000011110000;
		13'd3050: color_o = 12'b000011110000;
		13'd3051: color_o = 12'b000011110000;
		13'd3052: color_o = 12'b000011110000;
		13'd3053: color_o = 12'b000011110000;
		13'd3054: color_o = 12'b000011110000;
		13'd3055: color_o = 12'b000011110000;
		13'd3056: color_o = 12'b000011110000;
		13'd3057: color_o = 12'b000011110000;
		13'd3058: color_o = 12'b000011110000;
		13'd3059: color_o = 12'b000011110000;
		13'd3060: color_o = 12'b000011110000;
		13'd3061: color_o = 12'b000011110000;
		13'd3062: color_o = 12'b000011110000;
		13'd3063: color_o = 12'b000011110000;
		13'd3064: color_o = 12'b000011110000;
		13'd3065: color_o = 12'b000011110000;
		13'd3066: color_o = 12'b000011110000;
		13'd3067: color_o = 12'b000011110000;
		13'd3068: color_o = 12'b000011110000;
		13'd3069: color_o = 12'b000011110000;
		13'd3070: color_o = 12'b000011110000;
		13'd3071: color_o = 12'b000011110000;
		13'd3072: color_o = 12'b000011110000;
		13'd3073: color_o = 12'b000011110000;
		13'd3074: color_o = 12'b000011110000;
		13'd3075: color_o = 12'b000011110000;
		13'd3076: color_o = 12'b000011110000;
		13'd3077: color_o = 12'b000011110000;
		13'd3078: color_o = 12'b000011110000;
		13'd3079: color_o = 12'b000011110000;
		13'd3080: color_o = 12'b000011110000;
		13'd3081: color_o = 12'b000011110000;
		13'd3082: color_o = 12'b000000000000;
		13'd3083: color_o = 12'b000000000000;
		13'd3084: color_o = 12'b000000000000;
		13'd3085: color_o = 12'b000000000000;
		13'd3086: color_o = 12'b100000000000;
		13'd3087: color_o = 12'b100000000000;
		13'd3088: color_o = 12'b100000000000;
		13'd3089: color_o = 12'b100000000000;
		13'd3090: color_o = 12'b100000000000;
		13'd3091: color_o = 12'b100000000000;
		13'd3092: color_o = 12'b100000000000;
		13'd3093: color_o = 12'b100000000000;
		13'd3094: color_o = 12'b100000000000;
		13'd3095: color_o = 12'b100000000000;
		13'd3096: color_o = 12'b100000000000;
		13'd3097: color_o = 12'b100000000000;
		13'd3098: color_o = 12'b011000000000;
		13'd3099: color_o = 12'b011000000000;
		13'd3100: color_o = 12'b011000000000;
		13'd3101: color_o = 12'b011000000000;
		13'd3102: color_o = 12'b011000000000;
		13'd3103: color_o = 12'b000011110000;
		13'd3104: color_o = 12'b000011110000;
		13'd3105: color_o = 12'b000011110000;
		13'd3106: color_o = 12'b000011110000;
		13'd3107: color_o = 12'b000011110000;
		13'd3108: color_o = 12'b000011110000;
		13'd3109: color_o = 12'b000011110000;
		13'd3110: color_o = 12'b000011110000;
		13'd3111: color_o = 12'b000011110000;
		13'd3112: color_o = 12'b000011110000;
		13'd3113: color_o = 12'b000011110000;
		13'd3114: color_o = 12'b000011110000;
		13'd3115: color_o = 12'b000011110000;
		13'd3116: color_o = 12'b000011110000;
		13'd3117: color_o = 12'b000011110000;
		13'd3118: color_o = 12'b000011110000;
		13'd3119: color_o = 12'b000011110000;
		13'd3120: color_o = 12'b000011110000;
		13'd3121: color_o = 12'b000011110000;
		13'd3122: color_o = 12'b000011110000;
		13'd3123: color_o = 12'b000011110000;
		13'd3124: color_o = 12'b000011110000;
		13'd3125: color_o = 12'b000011110000;
		13'd3126: color_o = 12'b000011110000;
		13'd3127: color_o = 12'b000011110000;
		13'd3128: color_o = 12'b000011110000;
		13'd3129: color_o = 12'b000011110000;
		13'd3130: color_o = 12'b000011110000;
		13'd3131: color_o = 12'b000011110000;
		13'd3132: color_o = 12'b000011110000;
		13'd3133: color_o = 12'b000011110000;
		13'd3134: color_o = 12'b000011110000;
		13'd3135: color_o = 12'b000011110000;
		13'd3136: color_o = 12'b000011110000;
		13'd3137: color_o = 12'b000011110000;
		13'd3138: color_o = 12'b000011110000;
		13'd3139: color_o = 12'b000011110000;
		13'd3140: color_o = 12'b000011110000;
		13'd3141: color_o = 12'b000011110000;
		13'd3142: color_o = 12'b000011110000;
		13'd3143: color_o = 12'b000011110000;
		13'd3144: color_o = 12'b000011110000;
		13'd3145: color_o = 12'b000000000000;
		13'd3146: color_o = 12'b000000000000;
		13'd3147: color_o = 12'b100001000000;
		13'd3148: color_o = 12'b000000000000;
		13'd3149: color_o = 12'b000000000000;
		13'd3150: color_o = 12'b000000000000;
		13'd3151: color_o = 12'b000000000000;
		13'd3152: color_o = 12'b100000000000;
		13'd3153: color_o = 12'b100000000000;
		13'd3154: color_o = 12'b100000000000;
		13'd3155: color_o = 12'b100000000000;
		13'd3156: color_o = 12'b100000000000;
		13'd3157: color_o = 12'b100000000000;
		13'd3158: color_o = 12'b011000000000;
		13'd3159: color_o = 12'b011000000000;
		13'd3160: color_o = 12'b011000000000;
		13'd3161: color_o = 12'b100000000000;
		13'd3162: color_o = 12'b100000000000;
		13'd3163: color_o = 12'b100000000000;
		13'd3164: color_o = 12'b011000000000;
		13'd3165: color_o = 12'b011000000000;
		13'd3166: color_o = 12'b011000000000;
		13'd3167: color_o = 12'b011000000000;
		13'd3168: color_o = 12'b000011110000;
		13'd3169: color_o = 12'b000011110000;
		13'd3170: color_o = 12'b000011110000;
		13'd3171: color_o = 12'b000011110000;
		13'd3172: color_o = 12'b000011110000;
		13'd3173: color_o = 12'b000011110000;
		13'd3174: color_o = 12'b000011110000;
		13'd3175: color_o = 12'b000011110000;
		13'd3176: color_o = 12'b000011110000;
		13'd3177: color_o = 12'b000011110000;
		13'd3178: color_o = 12'b000011110000;
		13'd3179: color_o = 12'b000011110000;
		13'd3180: color_o = 12'b000011110000;
		13'd3181: color_o = 12'b000011110000;
		13'd3182: color_o = 12'b000011110000;
		13'd3183: color_o = 12'b000011110000;
		13'd3184: color_o = 12'b000011110000;
		13'd3185: color_o = 12'b000011110000;
		13'd3186: color_o = 12'b000011110000;
		13'd3187: color_o = 12'b000011110000;
		13'd3188: color_o = 12'b000011110000;
		13'd3189: color_o = 12'b000011110000;
		13'd3190: color_o = 12'b000011110000;
		13'd3191: color_o = 12'b000011110000;
		13'd3192: color_o = 12'b000011110000;
		13'd3193: color_o = 12'b000011110000;
		13'd3194: color_o = 12'b000011110000;
		13'd3195: color_o = 12'b000011110000;
		13'd3196: color_o = 12'b000011110000;
		13'd3197: color_o = 12'b000011110000;
		13'd3198: color_o = 12'b000011110000;
		13'd3199: color_o = 12'b000011110000;
		13'd3200: color_o = 12'b000011110000;
		13'd3201: color_o = 12'b000011110000;
		13'd3202: color_o = 12'b000011110000;
		13'd3203: color_o = 12'b000011110000;
		13'd3204: color_o = 12'b000011110000;
		13'd3205: color_o = 12'b000011110000;
		13'd3206: color_o = 12'b000011110000;
		13'd3207: color_o = 12'b000011110000;
		13'd3208: color_o = 12'b100001000000;
		13'd3209: color_o = 12'b100001000000;
		13'd3210: color_o = 12'b100001000000;
		13'd3211: color_o = 12'b000000000000;
		13'd3212: color_o = 12'b000000000000;
		13'd3213: color_o = 12'b100000000001;
		13'd3214: color_o = 12'b100000000001;
		13'd3215: color_o = 12'b100000000001;
		13'd3216: color_o = 12'b100000000001;
		13'd3217: color_o = 12'b000000000000;
		13'd3218: color_o = 12'b000000000000;
		13'd3219: color_o = 12'b000000000000;
		13'd3220: color_o = 12'b100000000000;
		13'd3221: color_o = 12'b100000000000;
		13'd3222: color_o = 12'b100000000000;
		13'd3223: color_o = 12'b100000000000;
		13'd3224: color_o = 12'b100000000000;
		13'd3225: color_o = 12'b100000000000;
		13'd3226: color_o = 12'b011000000000;
		13'd3227: color_o = 12'b011000000000;
		13'd3228: color_o = 12'b011000000000;
		13'd3229: color_o = 12'b011000000000;
		13'd3230: color_o = 12'b100000000000;
		13'd3231: color_o = 12'b100000000000;
		13'd3232: color_o = 12'b100000000000;
		13'd3233: color_o = 12'b000011110000;
		13'd3234: color_o = 12'b000011110000;
		13'd3235: color_o = 12'b000011110000;
		13'd3236: color_o = 12'b000011110000;
		13'd3237: color_o = 12'b000011110000;
		13'd3238: color_o = 12'b000011110000;
		13'd3239: color_o = 12'b000011110000;
		13'd3240: color_o = 12'b000011110000;
		13'd3241: color_o = 12'b000011110000;
		13'd3242: color_o = 12'b000011110000;
		13'd3243: color_o = 12'b000011110000;
		13'd3244: color_o = 12'b000011110000;
		13'd3245: color_o = 12'b000011110000;
		13'd3246: color_o = 12'b000011110000;
		13'd3247: color_o = 12'b000011110000;
		13'd3248: color_o = 12'b000011110000;
		13'd3249: color_o = 12'b000011110000;
		13'd3250: color_o = 12'b000011110000;
		13'd3251: color_o = 12'b000011110000;
		13'd3252: color_o = 12'b000011110000;
		13'd3253: color_o = 12'b000011110000;
		13'd3254: color_o = 12'b000011110000;
		13'd3255: color_o = 12'b000011110000;
		13'd3256: color_o = 12'b000011110000;
		13'd3257: color_o = 12'b000011110000;
		13'd3258: color_o = 12'b000011110000;
		13'd3259: color_o = 12'b000011110000;
		13'd3260: color_o = 12'b000011110000;
		13'd3261: color_o = 12'b000011110000;
		13'd3262: color_o = 12'b000011110000;
		13'd3263: color_o = 12'b000011110000;
		13'd3264: color_o = 12'b000011110000;
		13'd3265: color_o = 12'b000011110000;
		13'd3266: color_o = 12'b000011110000;
		13'd3267: color_o = 12'b000011110000;
		13'd3268: color_o = 12'b000011110000;
		13'd3269: color_o = 12'b000011110000;
		13'd3270: color_o = 12'b000011110000;
		13'd3271: color_o = 12'b000011110000;
		13'd3272: color_o = 12'b100001000000;
		13'd3273: color_o = 12'b100001000000;
		13'd3274: color_o = 12'b000000000000;
		13'd3275: color_o = 12'b000000000000;
		13'd3276: color_o = 12'b100000000001;
		13'd3277: color_o = 12'b100000000001;
		13'd3278: color_o = 12'b100000000001;
		13'd3279: color_o = 12'b100000000001;
		13'd3280: color_o = 12'b100000000001;
		13'd3281: color_o = 12'b100000000001;
		13'd3282: color_o = 12'b100000000001;
		13'd3283: color_o = 12'b000000000000;
		13'd3284: color_o = 12'b000000000000;
		13'd3285: color_o = 12'b000000000000;
		13'd3286: color_o = 12'b000000000000;
		13'd3287: color_o = 12'b000000000000;
		13'd3288: color_o = 12'b000000000000;
		13'd3289: color_o = 12'b100000000000;
		13'd3290: color_o = 12'b100000000000;
		13'd3291: color_o = 12'b100000000000;
		13'd3292: color_o = 12'b100000000000;
		13'd3293: color_o = 12'b100000000000;
		13'd3294: color_o = 12'b100000000000;
		13'd3295: color_o = 12'b100000000000;
		13'd3296: color_o = 12'b100000000000;
		13'd3297: color_o = 12'b000011110000;
		13'd3298: color_o = 12'b000011110000;
		13'd3299: color_o = 12'b000011110000;
		13'd3300: color_o = 12'b000011110000;
		13'd3301: color_o = 12'b000011110000;
		13'd3302: color_o = 12'b000011110000;
		13'd3303: color_o = 12'b000011110000;
		13'd3304: color_o = 12'b000011110000;
		13'd3305: color_o = 12'b000011110000;
		13'd3306: color_o = 12'b000011110000;
		13'd3307: color_o = 12'b000011110000;
		13'd3308: color_o = 12'b000011110000;
		13'd3309: color_o = 12'b000011110000;
		13'd3310: color_o = 12'b000011110000;
		13'd3311: color_o = 12'b000011110000;
		13'd3312: color_o = 12'b000011110000;
		13'd3313: color_o = 12'b000011110000;
		13'd3314: color_o = 12'b000011110000;
		13'd3315: color_o = 12'b000011110000;
		13'd3316: color_o = 12'b000011110000;
		13'd3317: color_o = 12'b000011110000;
		13'd3318: color_o = 12'b000011110000;
		13'd3319: color_o = 12'b000011110000;
		13'd3320: color_o = 12'b000011110000;
		13'd3321: color_o = 12'b000011110000;
		13'd3322: color_o = 12'b000011110000;
		13'd3323: color_o = 12'b000011110000;
		13'd3324: color_o = 12'b000011110000;
		13'd3325: color_o = 12'b000011110000;
		13'd3326: color_o = 12'b000011110000;
		13'd3327: color_o = 12'b000011110000;
		13'd3328: color_o = 12'b000011110000;
		13'd3329: color_o = 12'b000011110000;
		13'd3330: color_o = 12'b000011110000;
		13'd3331: color_o = 12'b000011110000;
		13'd3332: color_o = 12'b000011110000;
		13'd3333: color_o = 12'b000011110000;
		13'd3334: color_o = 12'b000011110000;
		13'd3335: color_o = 12'b000011110000;
		13'd3336: color_o = 12'b000000000000;
		13'd3337: color_o = 12'b000000000000;
		13'd3338: color_o = 12'b000000000000;
		13'd3339: color_o = 12'b100000000001;
		13'd3340: color_o = 12'b100000000001;
		13'd3341: color_o = 12'b100000000001;
		13'd3342: color_o = 12'b100000000001;
		13'd3343: color_o = 12'b100000000001;
		13'd3344: color_o = 12'b100000000001;
		13'd3345: color_o = 12'b000000000000;
		13'd3346: color_o = 12'b000000000000;
		13'd3347: color_o = 12'b000000000000;
		13'd3348: color_o = 12'b000000000000;
		13'd3349: color_o = 12'b000000000000;
		13'd3350: color_o = 12'b100000000001;
		13'd3351: color_o = 12'b100000000001;
		13'd3352: color_o = 12'b000000000000;
		13'd3353: color_o = 12'b000000000000;
		13'd3354: color_o = 12'b100000000000;
		13'd3355: color_o = 12'b100000000000;
		13'd3356: color_o = 12'b100000000000;
		13'd3357: color_o = 12'b100000000000;
		13'd3358: color_o = 12'b100000000000;
		13'd3359: color_o = 12'b100000000000;
		13'd3360: color_o = 12'b100000000000;
		13'd3361: color_o = 12'b000011110000;
		13'd3362: color_o = 12'b000011110000;
		13'd3363: color_o = 12'b000011110000;
		13'd3364: color_o = 12'b000011110000;
		13'd3365: color_o = 12'b000011110000;
		13'd3366: color_o = 12'b000011110000;
		13'd3367: color_o = 12'b000011110000;
		13'd3368: color_o = 12'b000011110000;
		13'd3369: color_o = 12'b000011110000;
		13'd3370: color_o = 12'b000011110000;
		13'd3371: color_o = 12'b000011110000;
		13'd3372: color_o = 12'b000011110000;
		13'd3373: color_o = 12'b000011110000;
		13'd3374: color_o = 12'b000011110000;
		13'd3375: color_o = 12'b000011110000;
		13'd3376: color_o = 12'b000011110000;
		13'd3377: color_o = 12'b000011110000;
		13'd3378: color_o = 12'b000011110000;
		13'd3379: color_o = 12'b000011110000;
		13'd3380: color_o = 12'b000011110000;
		13'd3381: color_o = 12'b000011110000;
		13'd3382: color_o = 12'b000011110000;
		13'd3383: color_o = 12'b000011110000;
		13'd3384: color_o = 12'b000011110000;
		13'd3385: color_o = 12'b000011110000;
		13'd3386: color_o = 12'b000011110000;
		13'd3387: color_o = 12'b000011110000;
		13'd3388: color_o = 12'b000011110000;
		13'd3389: color_o = 12'b000011110000;
		13'd3390: color_o = 12'b000011110000;
		13'd3391: color_o = 12'b000011110000;
		13'd3392: color_o = 12'b000011110000;
		13'd3393: color_o = 12'b000011110000;
		13'd3394: color_o = 12'b000011110000;
		13'd3395: color_o = 12'b000011110000;
		13'd3396: color_o = 12'b000011110000;
		13'd3397: color_o = 12'b000011110000;
		13'd3398: color_o = 12'b000011110000;
		13'd3399: color_o = 12'b000011110000;
		13'd3400: color_o = 12'b000000000000;
		13'd3401: color_o = 12'b000000000000;
		13'd3402: color_o = 12'b100000000001;
		13'd3403: color_o = 12'b100000000001;
		13'd3404: color_o = 12'b100000000001;
		13'd3405: color_o = 12'b000000000000;
		13'd3406: color_o = 12'b000000000000;
		13'd3407: color_o = 12'b000000000000;
		13'd3408: color_o = 12'b000000000000;
		13'd3409: color_o = 12'b000000000000;
		13'd3410: color_o = 12'b100000000001;
		13'd3411: color_o = 12'b100000000001;
		13'd3412: color_o = 12'b100000000001;
		13'd3413: color_o = 12'b100000000001;
		13'd3414: color_o = 12'b100000000001;
		13'd3415: color_o = 12'b100000000001;
		13'd3416: color_o = 12'b100000000001;
		13'd3417: color_o = 12'b000000000000;
		13'd3418: color_o = 12'b000000000000;
		13'd3419: color_o = 12'b000000000000;
		13'd3420: color_o = 12'b000000000000;
		13'd3421: color_o = 12'b000000000000;
		13'd3422: color_o = 12'b000000000000;
		13'd3423: color_o = 12'b000000000000;
		13'd3424: color_o = 12'b000000000000;
		13'd3425: color_o = 12'b111000010010;
		13'd3426: color_o = 12'b000011110000;
		13'd3427: color_o = 12'b000011110000;
		13'd3428: color_o = 12'b000011110000;
		13'd3429: color_o = 12'b000011110000;
		13'd3430: color_o = 12'b000011110000;
		13'd3431: color_o = 12'b000011110000;
		13'd3432: color_o = 12'b000011110000;
		13'd3433: color_o = 12'b000011110000;
		13'd3434: color_o = 12'b000011110000;
		13'd3435: color_o = 12'b000011110000;
		13'd3436: color_o = 12'b000011110000;
		13'd3437: color_o = 12'b000011110000;
		13'd3438: color_o = 12'b000011110000;
		13'd3439: color_o = 12'b000011110000;
		13'd3440: color_o = 12'b000011110000;
		13'd3441: color_o = 12'b000011110000;
		13'd3442: color_o = 12'b000011110000;
		13'd3443: color_o = 12'b000011110000;
		13'd3444: color_o = 12'b000011110000;
		13'd3445: color_o = 12'b000011110000;
		13'd3446: color_o = 12'b000011110000;
		13'd3447: color_o = 12'b000011110000;
		13'd3448: color_o = 12'b000011110000;
		13'd3449: color_o = 12'b000011110000;
		13'd3450: color_o = 12'b000011110000;
		13'd3451: color_o = 12'b000011110000;
		13'd3452: color_o = 12'b000011110000;
		13'd3453: color_o = 12'b000011110000;
		13'd3454: color_o = 12'b000011110000;
		13'd3455: color_o = 12'b000011110000;
		13'd3456: color_o = 12'b000011110000;
		13'd3457: color_o = 12'b000011110000;
		13'd3458: color_o = 12'b000011110000;
		13'd3459: color_o = 12'b000011110000;
		13'd3460: color_o = 12'b000011110000;
		13'd3461: color_o = 12'b000011110000;
		13'd3462: color_o = 12'b000011110000;
		13'd3463: color_o = 12'b000011110000;
		13'd3464: color_o = 12'b000000000000;
		13'd3465: color_o = 12'b000000000000;
		13'd3466: color_o = 12'b100000000001;
		13'd3467: color_o = 12'b000000000000;
		13'd3468: color_o = 12'b000000000000;
		13'd3469: color_o = 12'b000000000000;
		13'd3470: color_o = 12'b100001000000;
		13'd3471: color_o = 12'b100001000000;
		13'd3472: color_o = 12'b000000000000;
		13'd3473: color_o = 12'b100000000001;
		13'd3474: color_o = 12'b100000000001;
		13'd3475: color_o = 12'b100000000001;
		13'd3476: color_o = 12'b000000000000;
		13'd3477: color_o = 12'b000000000000;
		13'd3478: color_o = 12'b000000000000;
		13'd3479: color_o = 12'b000000000000;
		13'd3480: color_o = 12'b000000000000;
		13'd3481: color_o = 12'b111000010010;
		13'd3482: color_o = 12'b111000010010;
		13'd3483: color_o = 12'b111000010010;
		13'd3484: color_o = 12'b111000010010;
		13'd3485: color_o = 12'b111000010010;
		13'd3486: color_o = 12'b111000010010;
		13'd3487: color_o = 12'b111000010010;
		13'd3488: color_o = 12'b111000010010;
		13'd3489: color_o = 12'b111000010010;
		13'd3490: color_o = 12'b111000010010;
		13'd3491: color_o = 12'b000011110000;
		13'd3492: color_o = 12'b000011110000;
		13'd3493: color_o = 12'b000011110000;
		13'd3494: color_o = 12'b000011110000;
		13'd3495: color_o = 12'b000011110000;
		13'd3496: color_o = 12'b000011110000;
		13'd3497: color_o = 12'b000011110000;
		13'd3498: color_o = 12'b000011110000;
		13'd3499: color_o = 12'b000011110000;
		13'd3500: color_o = 12'b000011110000;
		13'd3501: color_o = 12'b000011110000;
		13'd3502: color_o = 12'b000011110000;
		13'd3503: color_o = 12'b000011110000;
		13'd3504: color_o = 12'b000011110000;
		13'd3505: color_o = 12'b000011110000;
		13'd3506: color_o = 12'b000011110000;
		13'd3507: color_o = 12'b000011110000;
		13'd3508: color_o = 12'b000011110000;
		13'd3509: color_o = 12'b000011110000;
		13'd3510: color_o = 12'b000011110000;
		13'd3511: color_o = 12'b000011110000;
		13'd3512: color_o = 12'b000011110000;
		13'd3513: color_o = 12'b000011110000;
		13'd3514: color_o = 12'b000011110000;
		13'd3515: color_o = 12'b000011110000;
		13'd3516: color_o = 12'b000011110000;
		13'd3517: color_o = 12'b000011110000;
		13'd3518: color_o = 12'b000011110000;
		13'd3519: color_o = 12'b000011110000;
		13'd3520: color_o = 12'b000011110000;
		13'd3521: color_o = 12'b000011110000;
		13'd3522: color_o = 12'b000011110000;
		13'd3523: color_o = 12'b000011110000;
		13'd3524: color_o = 12'b000011110000;
		13'd3525: color_o = 12'b000011110000;
		13'd3526: color_o = 12'b000011110000;
		13'd3527: color_o = 12'b000011110000;
		13'd3528: color_o = 12'b000000000000;
		13'd3529: color_o = 12'b000000000000;
		13'd3530: color_o = 12'b100000000001;
		13'd3531: color_o = 12'b000000000000;
		13'd3532: color_o = 12'b100001000000;
		13'd3533: color_o = 12'b100001000000;
		13'd3534: color_o = 12'b100001000000;
		13'd3535: color_o = 12'b100001000000;
		13'd3536: color_o = 12'b000000000000;
		13'd3537: color_o = 12'b100000000001;
		13'd3538: color_o = 12'b100000000001;
		13'd3539: color_o = 12'b000000000000;
		13'd3540: color_o = 12'b000000000000;
		13'd3541: color_o = 12'b000000000000;
		13'd3542: color_o = 12'b000000000000;
		13'd3543: color_o = 12'b000000000000;
		13'd3544: color_o = 12'b000000000000;
		13'd3545: color_o = 12'b000000000000;
		13'd3546: color_o = 12'b000000000000;
		13'd3547: color_o = 12'b000000000000;
		13'd3548: color_o = 12'b000000000000;
		13'd3549: color_o = 12'b000000000000;
		13'd3550: color_o = 12'b000000000000;
		13'd3551: color_o = 12'b000000000000;
		13'd3552: color_o = 12'b000000000000;
		13'd3553: color_o = 12'b000011110000;
		13'd3554: color_o = 12'b000011110000;
		13'd3555: color_o = 12'b000011110000;
		13'd3556: color_o = 12'b000011110000;
		13'd3557: color_o = 12'b000011110000;
		13'd3558: color_o = 12'b000011110000;
		13'd3559: color_o = 12'b000011110000;
		13'd3560: color_o = 12'b000011110000;
		13'd3561: color_o = 12'b000011110000;
		13'd3562: color_o = 12'b000011110000;
		13'd3563: color_o = 12'b000011110000;
		13'd3564: color_o = 12'b000011110000;
		13'd3565: color_o = 12'b000011110000;
		13'd3566: color_o = 12'b000011110000;
		13'd3567: color_o = 12'b000011110000;
		13'd3568: color_o = 12'b000011110000;
		13'd3569: color_o = 12'b000011110000;
		13'd3570: color_o = 12'b000011110000;
		13'd3571: color_o = 12'b000011110000;
		13'd3572: color_o = 12'b000011110000;
		13'd3573: color_o = 12'b000011110000;
		13'd3574: color_o = 12'b000011110000;
		13'd3575: color_o = 12'b000011110000;
		13'd3576: color_o = 12'b000011110000;
		13'd3577: color_o = 12'b000011110000;
		13'd3578: color_o = 12'b000011110000;
		13'd3579: color_o = 12'b000011110000;
		13'd3580: color_o = 12'b000011110000;
		13'd3581: color_o = 12'b000011110000;
		13'd3582: color_o = 12'b000011110000;
		13'd3583: color_o = 12'b000011110000;
		13'd3584: color_o = 12'b000011110000;
		13'd3585: color_o = 12'b000011110000;
		13'd3586: color_o = 12'b000011110000;
		13'd3587: color_o = 12'b000011110000;
		13'd3588: color_o = 12'b000011110000;
		13'd3589: color_o = 12'b000011110000;
		13'd3590: color_o = 12'b000011110000;
		13'd3591: color_o = 12'b000011110000;
		13'd3592: color_o = 12'b000000000000;
		13'd3593: color_o = 12'b000000000000;
		13'd3594: color_o = 12'b100000000001;
		13'd3595: color_o = 12'b000000000000;
		13'd3596: color_o = 12'b100001000000;
		13'd3597: color_o = 12'b100001000000;
		13'd3598: color_o = 12'b100001000000;
		13'd3599: color_o = 12'b100001000000;
		13'd3600: color_o = 12'b000000000000;
		13'd3601: color_o = 12'b100000000001;
		13'd3602: color_o = 12'b100000000001;
		13'd3603: color_o = 12'b000000000000;
		13'd3604: color_o = 12'b000000000000;
		13'd3605: color_o = 12'b000000000000;
		13'd3606: color_o = 12'b000000000000;
		13'd3607: color_o = 12'b000000000000;
		13'd3608: color_o = 12'b000000000000;
		13'd3609: color_o = 12'b000000000000;
		13'd3610: color_o = 12'b110011001100;
		13'd3611: color_o = 12'b110011001100;
		13'd3612: color_o = 12'b110011001100;
		13'd3613: color_o = 12'b000000000000;
		13'd3614: color_o = 12'b000000000000;
		13'd3615: color_o = 12'b000000000000;
		13'd3616: color_o = 12'b000000000000;
		13'd3617: color_o = 12'b000011110000;
		13'd3618: color_o = 12'b000011110000;
		13'd3619: color_o = 12'b000011110000;
		13'd3620: color_o = 12'b000011110000;
		13'd3621: color_o = 12'b000011110000;
		13'd3622: color_o = 12'b000011110000;
		13'd3623: color_o = 12'b000011110000;
		13'd3624: color_o = 12'b000011110000;
		13'd3625: color_o = 12'b000011110000;
		13'd3626: color_o = 12'b000011110000;
		13'd3627: color_o = 12'b000011110000;
		13'd3628: color_o = 12'b000011110000;
		13'd3629: color_o = 12'b000011110000;
		13'd3630: color_o = 12'b000011110000;
		13'd3631: color_o = 12'b000011110000;
		13'd3632: color_o = 12'b000011110000;
		13'd3633: color_o = 12'b000011110000;
		13'd3634: color_o = 12'b000011110000;
		13'd3635: color_o = 12'b000011110000;
		13'd3636: color_o = 12'b000011110000;
		13'd3637: color_o = 12'b000011110000;
		13'd3638: color_o = 12'b000011110000;
		13'd3639: color_o = 12'b000011110000;
		13'd3640: color_o = 12'b000011110000;
		13'd3641: color_o = 12'b000011110000;
		13'd3642: color_o = 12'b000011110000;
		13'd3643: color_o = 12'b000011110000;
		13'd3644: color_o = 12'b000011110000;
		13'd3645: color_o = 12'b000011110000;
		13'd3646: color_o = 12'b000011110000;
		13'd3647: color_o = 12'b000011110000;
		13'd3648: color_o = 12'b000011110000;
		13'd3649: color_o = 12'b000011110000;
		13'd3650: color_o = 12'b000011110000;
		13'd3651: color_o = 12'b000011110000;
		13'd3652: color_o = 12'b000011110000;
		13'd3653: color_o = 12'b000011110000;
		13'd3654: color_o = 12'b000011110000;
		13'd3655: color_o = 12'b000011110000;
		13'd3656: color_o = 12'b000000000000;
		13'd3657: color_o = 12'b100000000001;
		13'd3658: color_o = 12'b100000000001;
		13'd3659: color_o = 12'b000000000000;
		13'd3660: color_o = 12'b100001000000;
		13'd3661: color_o = 12'b100001000000;
		13'd3662: color_o = 12'b100001000000;
		13'd3663: color_o = 12'b100001000000;
		13'd3664: color_o = 12'b000000000000;
		13'd3665: color_o = 12'b100000000001;
		13'd3666: color_o = 12'b000000000000;
		13'd3667: color_o = 12'b000000000000;
		13'd3668: color_o = 12'b000000000000;
		13'd3669: color_o = 12'b000000000000;
		13'd3670: color_o = 12'b000000000000;
		13'd3671: color_o = 12'b000000000000;
		13'd3672: color_o = 12'b000000000000;
		13'd3673: color_o = 12'b000000000000;
		13'd3674: color_o = 12'b110011001100;
		13'd3675: color_o = 12'b110011001100;
		13'd3676: color_o = 12'b110011001100;
		13'd3677: color_o = 12'b000000000000;
		13'd3678: color_o = 12'b000000000000;
		13'd3679: color_o = 12'b000000000000;
		13'd3680: color_o = 12'b000000000000;
		13'd3681: color_o = 12'b000011110000;
		13'd3682: color_o = 12'b000011110000;
		13'd3683: color_o = 12'b000011110000;
		13'd3684: color_o = 12'b000011110000;
		13'd3685: color_o = 12'b000011110000;
		13'd3686: color_o = 12'b000011110000;
		13'd3687: color_o = 12'b000011110000;
		13'd3688: color_o = 12'b000011110000;
		13'd3689: color_o = 12'b000011110000;
		13'd3690: color_o = 12'b000011110000;
		13'd3691: color_o = 12'b000011110000;
		13'd3692: color_o = 12'b000011110000;
		13'd3693: color_o = 12'b000011110000;
		13'd3694: color_o = 12'b000011110000;
		13'd3695: color_o = 12'b000011110000;
		13'd3696: color_o = 12'b000011110000;
		13'd3697: color_o = 12'b000011110000;
		13'd3698: color_o = 12'b000011110000;
		13'd3699: color_o = 12'b000011110000;
		13'd3700: color_o = 12'b000011110000;
		13'd3701: color_o = 12'b000011110000;
		13'd3702: color_o = 12'b000011110000;
		13'd3703: color_o = 12'b000011110000;
		13'd3704: color_o = 12'b000011110000;
		13'd3705: color_o = 12'b000011110000;
		13'd3706: color_o = 12'b000011110000;
		13'd3707: color_o = 12'b000011110000;
		13'd3708: color_o = 12'b000011110000;
		13'd3709: color_o = 12'b000011110000;
		13'd3710: color_o = 12'b000011110000;
		13'd3711: color_o = 12'b000011110000;
		13'd3712: color_o = 12'b000011110000;
		13'd3713: color_o = 12'b000011110000;
		13'd3714: color_o = 12'b000011110000;
		13'd3715: color_o = 12'b000011110000;
		13'd3716: color_o = 12'b000011110000;
		13'd3717: color_o = 12'b000011110000;
		13'd3718: color_o = 12'b000011110000;
		13'd3719: color_o = 12'b000011110000;
		13'd3720: color_o = 12'b000000000000;
		13'd3721: color_o = 12'b100000000001;
		13'd3722: color_o = 12'b100000000001;
		13'd3723: color_o = 12'b000000000000;
		13'd3724: color_o = 12'b000000000000;
		13'd3725: color_o = 12'b000000000000;
		13'd3726: color_o = 12'b100001000000;
		13'd3727: color_o = 12'b100001000000;
		13'd3728: color_o = 12'b000000000000;
		13'd3729: color_o = 12'b100000000001;
		13'd3730: color_o = 12'b100000000001;
		13'd3731: color_o = 12'b000000000000;
		13'd3732: color_o = 12'b000000000000;
		13'd3733: color_o = 12'b000000000000;
		13'd3734: color_o = 12'b000000000000;
		13'd3735: color_o = 12'b000000000000;
		13'd3736: color_o = 12'b000000000000;
		13'd3737: color_o = 12'b000000000000;
		13'd3738: color_o = 12'b000000000000;
		13'd3739: color_o = 12'b000000000000;
		13'd3740: color_o = 12'b110011001100;
		13'd3741: color_o = 12'b000000000000;
		13'd3742: color_o = 12'b000000000000;
		13'd3743: color_o = 12'b000000000000;
		13'd3744: color_o = 12'b000000000000;
		13'd3745: color_o = 12'b000011110000;
		13'd3746: color_o = 12'b000011110000;
		13'd3747: color_o = 12'b000011110000;
		13'd3748: color_o = 12'b000011110000;
		13'd3749: color_o = 12'b000011110000;
		13'd3750: color_o = 12'b000011110000;
		13'd3751: color_o = 12'b000011110000;
		13'd3752: color_o = 12'b000011110000;
		13'd3753: color_o = 12'b000011110000;
		13'd3754: color_o = 12'b000011110000;
		13'd3755: color_o = 12'b000011110000;
		13'd3756: color_o = 12'b000011110000;
		13'd3757: color_o = 12'b000011110000;
		13'd3758: color_o = 12'b000011110000;
		13'd3759: color_o = 12'b000011110000;
		13'd3760: color_o = 12'b000011110000;
		13'd3761: color_o = 12'b000011110000;
		13'd3762: color_o = 12'b000011110000;
		13'd3763: color_o = 12'b000011110000;
		13'd3764: color_o = 12'b000011110000;
		13'd3765: color_o = 12'b000011110000;
		13'd3766: color_o = 12'b000011110000;
		13'd3767: color_o = 12'b000011110000;
		13'd3768: color_o = 12'b000011110000;
		13'd3769: color_o = 12'b000011110000;
		13'd3770: color_o = 12'b000011110000;
		13'd3771: color_o = 12'b000011110000;
		13'd3772: color_o = 12'b000011110000;
		13'd3773: color_o = 12'b000011110000;
		13'd3774: color_o = 12'b000011110000;
		13'd3775: color_o = 12'b000011110000;
		13'd3776: color_o = 12'b000011110000;
		13'd3777: color_o = 12'b000011110000;
		13'd3778: color_o = 12'b000011110000;
		13'd3779: color_o = 12'b000011110000;
		13'd3780: color_o = 12'b000011110000;
		13'd3781: color_o = 12'b000011110000;
		13'd3782: color_o = 12'b000011110000;
		13'd3783: color_o = 12'b000011110000;
		13'd3784: color_o = 12'b100000000001;
		13'd3785: color_o = 12'b100000000001;
		13'd3786: color_o = 12'b100000000001;
		13'd3787: color_o = 12'b100000000001;
		13'd3788: color_o = 12'b000000000000;
		13'd3789: color_o = 12'b000000000000;
		13'd3790: color_o = 12'b000000000000;
		13'd3791: color_o = 12'b000000000000;
		13'd3792: color_o = 12'b000000000000;
		13'd3793: color_o = 12'b000000000000;
		13'd3794: color_o = 12'b100000000001;
		13'd3795: color_o = 12'b100000000001;
		13'd3796: color_o = 12'b000000000000;
		13'd3797: color_o = 12'b000000000000;
		13'd3798: color_o = 12'b000000000000;
		13'd3799: color_o = 12'b000000000000;
		13'd3800: color_o = 12'b000000000000;
		13'd3801: color_o = 12'b000000000000;
		13'd3802: color_o = 12'b000000000000;
		13'd3803: color_o = 12'b000000000000;
		13'd3804: color_o = 12'b000000000000;
		13'd3805: color_o = 12'b000000000000;
		13'd3806: color_o = 12'b000000000000;
		13'd3807: color_o = 12'b000000000000;
		13'd3808: color_o = 12'b000011110000;
		13'd3809: color_o = 12'b000011110000;
		13'd3810: color_o = 12'b000011110000;
		13'd3811: color_o = 12'b000011110000;
		13'd3812: color_o = 12'b000011110000;
		13'd3813: color_o = 12'b000011110000;
		13'd3814: color_o = 12'b000011110000;
		13'd3815: color_o = 12'b000011110000;
		13'd3816: color_o = 12'b000011110000;
		13'd3817: color_o = 12'b000011110000;
		13'd3818: color_o = 12'b000011110000;
		13'd3819: color_o = 12'b000011110000;
		13'd3820: color_o = 12'b000011110000;
		13'd3821: color_o = 12'b000011110000;
		13'd3822: color_o = 12'b000011110000;
		13'd3823: color_o = 12'b000011110000;
		13'd3824: color_o = 12'b000011110000;
		13'd3825: color_o = 12'b000011110000;
		13'd3826: color_o = 12'b000011110000;
		13'd3827: color_o = 12'b000011110000;
		13'd3828: color_o = 12'b000011110000;
		13'd3829: color_o = 12'b000011110000;
		13'd3830: color_o = 12'b000011110000;
		13'd3831: color_o = 12'b000011110000;
		13'd3832: color_o = 12'b000011110000;
		13'd3833: color_o = 12'b000011110000;
		13'd3834: color_o = 12'b000011110000;
		13'd3835: color_o = 12'b000011110000;
		13'd3836: color_o = 12'b000011110000;
		13'd3837: color_o = 12'b000011110000;
		13'd3838: color_o = 12'b000011110000;
		13'd3839: color_o = 12'b000011110000;
		13'd3840: color_o = 12'b000011110000;
		13'd3841: color_o = 12'b000011110000;
		13'd3842: color_o = 12'b000011110000;
		13'd3843: color_o = 12'b000011110000;
		13'd3844: color_o = 12'b000011110000;
		13'd3845: color_o = 12'b000011110000;
		13'd3846: color_o = 12'b000011110000;
		13'd3847: color_o = 12'b000011110000;
		13'd3848: color_o = 12'b100000000001;
		13'd3849: color_o = 12'b100000000001;
		13'd3850: color_o = 12'b000000000000;
		13'd3851: color_o = 12'b000000000000;
		13'd3852: color_o = 12'b111000010010;
		13'd3853: color_o = 12'b111000010010;
		13'd3854: color_o = 12'b000000000000;
		13'd3855: color_o = 12'b000000000000;
		13'd3856: color_o = 12'b000000000000;
		13'd3857: color_o = 12'b000000000000;
		13'd3858: color_o = 12'b000000000000;
		13'd3859: color_o = 12'b000000000000;
		13'd3860: color_o = 12'b100000000001;
		13'd3861: color_o = 12'b100000000001;
		13'd3862: color_o = 12'b100000000001;
		13'd3863: color_o = 12'b100000000001;
		13'd3864: color_o = 12'b100000000001;
		13'd3865: color_o = 12'b100000000001;
		13'd3866: color_o = 12'b100000000001;
		13'd3867: color_o = 12'b100000000001;
		13'd3868: color_o = 12'b100000000001;
		13'd3869: color_o = 12'b100000000001;
		13'd3870: color_o = 12'b100000000001;
		13'd3871: color_o = 12'b100000000001;
		13'd3872: color_o = 12'b000011110000;
		13'd3873: color_o = 12'b000011110000;
		13'd3874: color_o = 12'b000011110000;
		13'd3875: color_o = 12'b000011110000;
		13'd3876: color_o = 12'b000011110000;
		13'd3877: color_o = 12'b000011110000;
		13'd3878: color_o = 12'b000011110000;
		13'd3879: color_o = 12'b000011110000;
		13'd3880: color_o = 12'b000011110000;
		13'd3881: color_o = 12'b000011110000;
		13'd3882: color_o = 12'b000011110000;
		13'd3883: color_o = 12'b000011110000;
		13'd3884: color_o = 12'b000000000000;
		13'd3885: color_o = 12'b000000000000;
		13'd3886: color_o = 12'b000000000000;
		13'd3887: color_o = 12'b000011110000;
		13'd3888: color_o = 12'b000011110000;
		13'd3889: color_o = 12'b000011110000;
		13'd3890: color_o = 12'b000011110000;
		13'd3891: color_o = 12'b000011110000;
		13'd3892: color_o = 12'b000011110000;
		13'd3893: color_o = 12'b000011110000;
		13'd3894: color_o = 12'b000011110000;
		13'd3895: color_o = 12'b000011110000;
		13'd3896: color_o = 12'b000011110000;
		13'd3897: color_o = 12'b000011110000;
		13'd3898: color_o = 12'b000011110000;
		13'd3899: color_o = 12'b000011110000;
		13'd3900: color_o = 12'b000011110000;
		13'd3901: color_o = 12'b000011110000;
		13'd3902: color_o = 12'b000011110000;
		13'd3903: color_o = 12'b000011110000;
		13'd3904: color_o = 12'b000011110000;
		13'd3905: color_o = 12'b000011110000;
		13'd3906: color_o = 12'b000011110000;
		13'd3907: color_o = 12'b000011110000;
		13'd3908: color_o = 12'b000011110000;
		13'd3909: color_o = 12'b000011110000;
		13'd3910: color_o = 12'b000011110000;
		13'd3911: color_o = 12'b000000000000;
		13'd3912: color_o = 12'b000000000000;
		13'd3913: color_o = 12'b100000000001;
		13'd3914: color_o = 12'b000000000000;
		13'd3915: color_o = 12'b111000010010;
		13'd3916: color_o = 12'b111000010010;
		13'd3917: color_o = 12'b000000000000;
		13'd3918: color_o = 12'b000000000000;
		13'd3919: color_o = 12'b100000000001;
		13'd3920: color_o = 12'b000000000000;
		13'd3921: color_o = 12'b111000010010;
		13'd3922: color_o = 12'b111000010010;
		13'd3923: color_o = 12'b000000000000;
		13'd3924: color_o = 12'b000000000000;
		13'd3925: color_o = 12'b000000000000;
		13'd3926: color_o = 12'b000000000000;
		13'd3927: color_o = 12'b000000000000;
		13'd3928: color_o = 12'b000000000000;
		13'd3929: color_o = 12'b000000000000;
		13'd3930: color_o = 12'b000000000000;
		13'd3931: color_o = 12'b000000000000;
		13'd3932: color_o = 12'b000000000000;
		13'd3933: color_o = 12'b100000000001;
		13'd3934: color_o = 12'b100000000001;
		13'd3935: color_o = 12'b100000000001;
		13'd3936: color_o = 12'b100000000001;
		13'd3937: color_o = 12'b000011110000;
		13'd3938: color_o = 12'b000011110000;
		13'd3939: color_o = 12'b000011110000;
		13'd3940: color_o = 12'b000011110000;
		13'd3941: color_o = 12'b000011110000;
		13'd3942: color_o = 12'b000011110000;
		13'd3943: color_o = 12'b000011110000;
		13'd3944: color_o = 12'b000011110000;
		13'd3945: color_o = 12'b000000000000;
		13'd3946: color_o = 12'b000000000000;
		13'd3947: color_o = 12'b000000000000;
		13'd3948: color_o = 12'b010001000100;
		13'd3949: color_o = 12'b010001000100;
		13'd3950: color_o = 12'b010001000100;
		13'd3951: color_o = 12'b000011110000;
		13'd3952: color_o = 12'b000011110000;
		13'd3953: color_o = 12'b000011110000;
		13'd3954: color_o = 12'b000011110000;
		13'd3955: color_o = 12'b000011110000;
		13'd3956: color_o = 12'b000011110000;
		13'd3957: color_o = 12'b000011110000;
		13'd3958: color_o = 12'b000011110000;
		13'd3959: color_o = 12'b000011110000;
		13'd3960: color_o = 12'b000011110000;
		13'd3961: color_o = 12'b000011110000;
		13'd3962: color_o = 12'b000011110000;
		13'd3963: color_o = 12'b000011110000;
		13'd3964: color_o = 12'b000011110000;
		13'd3965: color_o = 12'b000011110000;
		13'd3966: color_o = 12'b000011110000;
		13'd3967: color_o = 12'b000011110000;
		13'd3968: color_o = 12'b000011110000;
		13'd3969: color_o = 12'b000011110000;
		13'd3970: color_o = 12'b000011110000;
		13'd3971: color_o = 12'b000011110000;
		13'd3972: color_o = 12'b000011110000;
		13'd3973: color_o = 12'b000011110000;
		13'd3974: color_o = 12'b000000000000;
		13'd3975: color_o = 12'b000000000000;
		13'd3976: color_o = 12'b000000000000;
		13'd3977: color_o = 12'b000000000000;
		13'd3978: color_o = 12'b000000000000;
		13'd3979: color_o = 12'b100000000001;
		13'd3980: color_o = 12'b100000000001;
		13'd3981: color_o = 12'b000000000000;
		13'd3982: color_o = 12'b100000000000;
		13'd3983: color_o = 12'b100000000000;
		13'd3984: color_o = 12'b000000000000;
		13'd3985: color_o = 12'b000000000000;
		13'd3986: color_o = 12'b111000010010;
		13'd3987: color_o = 12'b000000000000;
		13'd3988: color_o = 12'b000000000000;
		13'd3989: color_o = 12'b100000000001;
		13'd3990: color_o = 12'b100000000001;
		13'd3991: color_o = 12'b100000000001;
		13'd3992: color_o = 12'b000000000000;
		13'd3993: color_o = 12'b111000010010;
		13'd3994: color_o = 12'b111000010010;
		13'd3995: color_o = 12'b000000000000;
		13'd3996: color_o = 12'b000000000000;
		13'd3997: color_o = 12'b100000000001;
		13'd3998: color_o = 12'b100000000001;
		13'd3999: color_o = 12'b100000000001;
		13'd4000: color_o = 12'b100000000001;
		13'd4001: color_o = 12'b000011110000;
		13'd4002: color_o = 12'b000011110000;
		13'd4003: color_o = 12'b000011110000;
		13'd4004: color_o = 12'b000011110000;
		13'd4005: color_o = 12'b000011110000;
		13'd4006: color_o = 12'b000011110000;
		13'd4007: color_o = 12'b000000000000;
		13'd4008: color_o = 12'b000000000000;
		13'd4009: color_o = 12'b010001000100;
		13'd4010: color_o = 12'b010001000100;
		13'd4011: color_o = 12'b010001000100;
		13'd4012: color_o = 12'b011101110111;
		13'd4013: color_o = 12'b011101110111;
		13'd4014: color_o = 12'b011101110111;
		13'd4015: color_o = 12'b000000000000;
		13'd4016: color_o = 12'b010001000100;
		13'd4017: color_o = 12'b000011110000;
		13'd4018: color_o = 12'b000011110000;
		13'd4019: color_o = 12'b000011110000;
		13'd4020: color_o = 12'b000011110000;
		13'd4021: color_o = 12'b000011110000;
		13'd4022: color_o = 12'b000011110000;
		13'd4023: color_o = 12'b000011110000;
		13'd4024: color_o = 12'b000011110000;
		13'd4025: color_o = 12'b000011110000;
		13'd4026: color_o = 12'b000011110000;
		13'd4027: color_o = 12'b000011110000;
		13'd4028: color_o = 12'b000011110000;
		13'd4029: color_o = 12'b000011110000;
		13'd4030: color_o = 12'b000011110000;
		13'd4031: color_o = 12'b000011110000;
		13'd4032: color_o = 12'b000011110000;
		13'd4033: color_o = 12'b000011110000;
		13'd4034: color_o = 12'b000011110000;
		13'd4035: color_o = 12'b000011110000;
		13'd4036: color_o = 12'b000011110000;
		13'd4037: color_o = 12'b000000000000;
		13'd4038: color_o = 12'b000000000000;
		13'd4039: color_o = 12'b000000000000;
		13'd4040: color_o = 12'b000000000000;
		13'd4041: color_o = 12'b100000000000;
		13'd4042: color_o = 12'b000000000000;
		13'd4043: color_o = 12'b000000000000;
		13'd4044: color_o = 12'b100000000000;
		13'd4045: color_o = 12'b000000000000;
		13'd4046: color_o = 12'b000000000000;
		13'd4047: color_o = 12'b000000000000;
		13'd4048: color_o = 12'b000000000000;
		13'd4049: color_o = 12'b000000000000;
		13'd4050: color_o = 12'b000000000000;
		13'd4051: color_o = 12'b000000000000;
		13'd4052: color_o = 12'b000000000000;
		13'd4053: color_o = 12'b100000000000;
		13'd4054: color_o = 12'b100000000000;
		13'd4055: color_o = 12'b000000000000;
		13'd4056: color_o = 12'b111000010010;
		13'd4057: color_o = 12'b111000010010;
		13'd4058: color_o = 12'b111000010010;
		13'd4059: color_o = 12'b000000000000;
		13'd4060: color_o = 12'b100000000001;
		13'd4061: color_o = 12'b100000000001;
		13'd4062: color_o = 12'b100000000001;
		13'd4063: color_o = 12'b100000000001;
		13'd4064: color_o = 12'b000000000000;
		13'd4065: color_o = 12'b000011110000;
		13'd4066: color_o = 12'b000011110000;
		13'd4067: color_o = 12'b000011110000;
		13'd4068: color_o = 12'b000000000000;
		13'd4069: color_o = 12'b000000000000;
		13'd4070: color_o = 12'b000000000000;
		13'd4071: color_o = 12'b010001000100;
		13'd4072: color_o = 12'b010001000100;
		13'd4073: color_o = 12'b011101110111;
		13'd4074: color_o = 12'b011101110111;
		13'd4075: color_o = 12'b011101110111;
		13'd4076: color_o = 12'b000000000000;
		13'd4077: color_o = 12'b000000000000;
		13'd4078: color_o = 12'b000000000000;
		13'd4079: color_o = 12'b011101110111;
		13'd4080: color_o = 12'b010001000100;
		13'd4081: color_o = 12'b000011110000;
		13'd4082: color_o = 12'b000011110000;
		13'd4083: color_o = 12'b000011110000;
		13'd4084: color_o = 12'b000011110000;
		13'd4085: color_o = 12'b000011110000;
		13'd4086: color_o = 12'b000011110000;
		13'd4087: color_o = 12'b000011110000;
		13'd4088: color_o = 12'b000011110000;
		13'd4089: color_o = 12'b000011110000;
		13'd4090: color_o = 12'b000011110000;
		13'd4091: color_o = 12'b000011110000;
		13'd4092: color_o = 12'b000011110000;
		13'd4093: color_o = 12'b000011110000;
		13'd4094: color_o = 12'b000011110000;
		13'd4095: color_o = 12'b000011110000;
		13'd4096: color_o = 12'b000011110000;
		13'd4097: color_o = 12'b000011110000;
		13'd4098: color_o = 12'b000011110000;
		13'd4099: color_o = 12'b000011110000;
		13'd4100: color_o = 12'b000011110000;
		13'd4101: color_o = 12'b000000000000;
		13'd4102: color_o = 12'b100001000000;
		13'd4103: color_o = 12'b000000000000;
		13'd4104: color_o = 12'b000000000000;
		13'd4105: color_o = 12'b100000000001;
		13'd4106: color_o = 12'b100000000000;
		13'd4107: color_o = 12'b000000000000;
		13'd4108: color_o = 12'b000000000000;
		13'd4109: color_o = 12'b000000000000;
		13'd4110: color_o = 12'b100000000000;
		13'd4111: color_o = 12'b100000000000;
		13'd4112: color_o = 12'b100000000000;
		13'd4113: color_o = 12'b000000000000;
		13'd4114: color_o = 12'b000000000000;
		13'd4115: color_o = 12'b100000000000;
		13'd4116: color_o = 12'b000000000000;
		13'd4117: color_o = 12'b000000000000;
		13'd4118: color_o = 12'b000000000000;
		13'd4119: color_o = 12'b000000000000;
		13'd4120: color_o = 12'b000000000000;
		13'd4121: color_o = 12'b111000010010;
		13'd4122: color_o = 12'b111000010010;
		13'd4123: color_o = 12'b000000000000;
		13'd4124: color_o = 12'b000000000000;
		13'd4125: color_o = 12'b000000000000;
		13'd4126: color_o = 12'b000000000000;
		13'd4127: color_o = 12'b000000000000;
		13'd4128: color_o = 12'b000000000000;
		13'd4129: color_o = 12'b000011110000;
		13'd4130: color_o = 12'b000000000000;
		13'd4131: color_o = 12'b000000000000;
		13'd4132: color_o = 12'b010001000100;
		13'd4133: color_o = 12'b010001000100;
		13'd4134: color_o = 12'b010001000100;
		13'd4135: color_o = 12'b011101110111;
		13'd4136: color_o = 12'b011101110111;
		13'd4137: color_o = 12'b000000000000;
		13'd4138: color_o = 12'b000000000000;
		13'd4139: color_o = 12'b000000000000;
		13'd4140: color_o = 12'b011101110111;
		13'd4141: color_o = 12'b011101110111;
		13'd4142: color_o = 12'b011101110111;
		13'd4143: color_o = 12'b011101110111;
		13'd4144: color_o = 12'b011101110111;
		13'd4145: color_o = 12'b000011110000;
		13'd4146: color_o = 12'b000011110000;
		13'd4147: color_o = 12'b000011110000;
		13'd4148: color_o = 12'b000011110000;
		13'd4149: color_o = 12'b000011110000;
		13'd4150: color_o = 12'b000011110000;
		13'd4151: color_o = 12'b000011110000;
		13'd4152: color_o = 12'b000011110000;
		13'd4153: color_o = 12'b000011110000;
		13'd4154: color_o = 12'b000011110000;
		13'd4155: color_o = 12'b000011110000;
		13'd4156: color_o = 12'b000011110000;
		13'd4157: color_o = 12'b000011110000;
		13'd4158: color_o = 12'b000011110000;
		13'd4159: color_o = 12'b000011110000;
		13'd4160: color_o = 12'b000011110000;
		13'd4161: color_o = 12'b000011110000;
		13'd4162: color_o = 12'b000011110000;
		13'd4163: color_o = 12'b000011110000;
		13'd4164: color_o = 12'b000000000000;
		13'd4165: color_o = 12'b000000000000;
		13'd4166: color_o = 12'b100001000000;
		13'd4167: color_o = 12'b000000000000;
		13'd4168: color_o = 12'b000000000000;
		13'd4169: color_o = 12'b100000000001;
		13'd4170: color_o = 12'b100000000000;
		13'd4171: color_o = 12'b000000000000;
		13'd4172: color_o = 12'b000000000000;
		13'd4173: color_o = 12'b100000000000;
		13'd4174: color_o = 12'b100000000000;
		13'd4175: color_o = 12'b100000000000;
		13'd4176: color_o = 12'b100000000000;
		13'd4177: color_o = 12'b100000000000;
		13'd4178: color_o = 12'b100000000000;
		13'd4179: color_o = 12'b100000000000;
		13'd4180: color_o = 12'b000000000000;
		13'd4181: color_o = 12'b100000000000;
		13'd4182: color_o = 12'b100000000000;
		13'd4183: color_o = 12'b000000000000;
		13'd4184: color_o = 12'b000000000000;
		13'd4185: color_o = 12'b000000000000;
		13'd4186: color_o = 12'b000000000000;
		13'd4187: color_o = 12'b000000000000;
		13'd4188: color_o = 12'b000000000000;
		13'd4189: color_o = 12'b000011110000;
		13'd4190: color_o = 12'b000011110000;
		13'd4191: color_o = 12'b000011110000;
		13'd4192: color_o = 12'b000011110000;
		13'd4193: color_o = 12'b000011110000;
		13'd4194: color_o = 12'b010001000100;
		13'd4195: color_o = 12'b010001000100;
		13'd4196: color_o = 12'b011101110111;
		13'd4197: color_o = 12'b011101110111;
		13'd4198: color_o = 12'b011101110111;
		13'd4199: color_o = 12'b000000000000;
		13'd4200: color_o = 12'b000000000000;
		13'd4201: color_o = 12'b011110011011;
		13'd4202: color_o = 12'b011101110111;
		13'd4203: color_o = 12'b011101110111;
		13'd4204: color_o = 12'b011010001010;
		13'd4205: color_o = 12'b011110011011;
		13'd4206: color_o = 12'b011101110111;
		13'd4207: color_o = 12'b011110011011;
		13'd4208: color_o = 12'b011101110111;
		13'd4209: color_o = 12'b011101110111;
		13'd4210: color_o = 12'b010001000100;
		13'd4211: color_o = 12'b000011110000;
		13'd4212: color_o = 12'b000011110000;
		13'd4213: color_o = 12'b000011110000;
		13'd4214: color_o = 12'b000011110000;
		13'd4215: color_o = 12'b000011110000;
		13'd4216: color_o = 12'b000011110000;
		13'd4217: color_o = 12'b000011110000;
		13'd4218: color_o = 12'b000011110000;
		13'd4219: color_o = 12'b000011110000;
		13'd4220: color_o = 12'b000011110000;
		13'd4221: color_o = 12'b000011110000;
		13'd4222: color_o = 12'b000011110000;
		13'd4223: color_o = 12'b000011110000;
		13'd4224: color_o = 12'b000011110000;
		13'd4225: color_o = 12'b000011110000;
		13'd4226: color_o = 12'b000011110000;
		13'd4227: color_o = 12'b000011110000;
		13'd4228: color_o = 12'b000000000000;
		13'd4229: color_o = 12'b100000000001;
		13'd4230: color_o = 12'b000000000000;
		13'd4231: color_o = 12'b000000000000;
		13'd4232: color_o = 12'b000000000000;
		13'd4233: color_o = 12'b100000000001;
		13'd4234: color_o = 12'b100000000000;
		13'd4235: color_o = 12'b000000000000;
		13'd4236: color_o = 12'b100000000000;
		13'd4237: color_o = 12'b000000000000;
		13'd4238: color_o = 12'b100000000000;
		13'd4239: color_o = 12'b010000000000;
		13'd4240: color_o = 12'b100000000000;
		13'd4241: color_o = 12'b000000000000;
		13'd4242: color_o = 12'b100000000000;
		13'd4243: color_o = 12'b100000000000;
		13'd4244: color_o = 12'b100000000000;
		13'd4245: color_o = 12'b000000000000;
		13'd4246: color_o = 12'b000000000000;
		13'd4247: color_o = 12'b000000000000;
		13'd4248: color_o = 12'b000000000000;
		13'd4249: color_o = 12'b010000000000;
		13'd4250: color_o = 12'b010000000000;
		13'd4251: color_o = 12'b000000000000;
		13'd4252: color_o = 12'b000011110000;
		13'd4253: color_o = 12'b000011110000;
		13'd4254: color_o = 12'b000000000000;
		13'd4255: color_o = 12'b000000000000;
		13'd4256: color_o = 12'b011110011011;
		13'd4257: color_o = 12'b011101110111;
		13'd4258: color_o = 12'b011101110111;
		13'd4259: color_o = 12'b011101110111;
		13'd4260: color_o = 12'b000000000000;
		13'd4261: color_o = 12'b000000000000;
		13'd4262: color_o = 12'b000000000000;
		13'd4263: color_o = 12'b011101110111;
		13'd4264: color_o = 12'b011110011011;
		13'd4265: color_o = 12'b011101110111;
		13'd4266: color_o = 12'b011101110111;
		13'd4267: color_o = 12'b011110011011;
		13'd4268: color_o = 12'b000000000000;
		13'd4269: color_o = 12'b000000000000;
		13'd4270: color_o = 12'b000000000000;
		13'd4271: color_o = 12'b011110011011;
		13'd4272: color_o = 12'b011110011011;
		13'd4273: color_o = 12'b011101110111;
		13'd4274: color_o = 12'b000000000000;
		13'd4275: color_o = 12'b000000000000;
		13'd4276: color_o = 12'b000011110000;
		13'd4277: color_o = 12'b000011110000;
		13'd4278: color_o = 12'b000011110000;
		13'd4279: color_o = 12'b000011110000;
		13'd4280: color_o = 12'b000011110000;
		13'd4281: color_o = 12'b000011110000;
		13'd4282: color_o = 12'b000011110000;
		13'd4283: color_o = 12'b000011110000;
		13'd4284: color_o = 12'b000011110000;
		13'd4285: color_o = 12'b000011110000;
		13'd4286: color_o = 12'b000011110000;
		13'd4287: color_o = 12'b000011110000;
		13'd4288: color_o = 12'b000011110000;
		13'd4289: color_o = 12'b000011110000;
		13'd4290: color_o = 12'b000011110000;
		13'd4291: color_o = 12'b000011110000;
		13'd4292: color_o = 12'b000000000000;
		13'd4293: color_o = 12'b100000000001;
		13'd4294: color_o = 12'b000000000000;
		13'd4295: color_o = 12'b100000000000;
		13'd4296: color_o = 12'b000000000000;
		13'd4297: color_o = 12'b100000000001;
		13'd4298: color_o = 12'b100000000000;
		13'd4299: color_o = 12'b000000000000;
		13'd4300: color_o = 12'b100000000000;
		13'd4301: color_o = 12'b000000000000;
		13'd4302: color_o = 12'b000000000000;
		13'd4303: color_o = 12'b010000000000;
		13'd4304: color_o = 12'b010000000000;
		13'd4305: color_o = 12'b000000000000;
		13'd4306: color_o = 12'b100000000000;
		13'd4307: color_o = 12'b100000000000;
		13'd4308: color_o = 12'b100000000000;
		13'd4309: color_o = 12'b000000000000;
		13'd4310: color_o = 12'b100000000001;
		13'd4311: color_o = 12'b100000000000;
		13'd4312: color_o = 12'b100000000000;
		13'd4313: color_o = 12'b000000000000;
		13'd4314: color_o = 12'b010000000000;
		13'd4315: color_o = 12'b010000000000;
		13'd4316: color_o = 12'b010000000000;
		13'd4317: color_o = 12'b010000000000;
		13'd4318: color_o = 12'b011110011011;
		13'd4319: color_o = 12'b011110011011;
		13'd4320: color_o = 12'b011110011011;
		13'd4321: color_o = 12'b000000000000;
		13'd4322: color_o = 12'b000000000000;
		13'd4323: color_o = 12'b000000000000;
		13'd4324: color_o = 12'b011110011011;
		13'd4325: color_o = 12'b011101110111;
		13'd4326: color_o = 12'b011101110111;
		13'd4327: color_o = 12'b011110011011;
		13'd4328: color_o = 12'b011101110111;
		13'd4329: color_o = 12'b000000000000;
		13'd4330: color_o = 12'b000000000000;
		13'd4331: color_o = 12'b000000000000;
		13'd4332: color_o = 12'b000000000000;
		13'd4333: color_o = 12'b011101110111;
		13'd4334: color_o = 12'b011110011011;
		13'd4335: color_o = 12'b011101110111;
		13'd4336: color_o = 12'b011101110111;
		13'd4337: color_o = 12'b000000000000;
		13'd4338: color_o = 12'b000011110000;
		13'd4339: color_o = 12'b000011110000;
		13'd4340: color_o = 12'b000011110000;
		13'd4341: color_o = 12'b000011110000;
		13'd4342: color_o = 12'b000011110000;
		13'd4343: color_o = 12'b000011110000;
		13'd4344: color_o = 12'b000011110000;
		13'd4345: color_o = 12'b000011110000;
		13'd4346: color_o = 12'b000011110000;
		13'd4347: color_o = 12'b000011110000;
		13'd4348: color_o = 12'b000011110000;
		13'd4349: color_o = 12'b000011110000;
		13'd4350: color_o = 12'b000011110000;
		13'd4351: color_o = 12'b000011110000;
		13'd4352: color_o = 12'b000011110000;
		13'd4353: color_o = 12'b000011110000;
		13'd4354: color_o = 12'b000011110000;
		13'd4355: color_o = 12'b000000000000;
		13'd4356: color_o = 12'b000000000000;
		13'd4357: color_o = 12'b100000000001;
		13'd4358: color_o = 12'b000000000000;
		13'd4359: color_o = 12'b000000000000;
		13'd4360: color_o = 12'b000000000000;
		13'd4361: color_o = 12'b100000000001;
		13'd4362: color_o = 12'b000000000000;
		13'd4363: color_o = 12'b100000000000;
		13'd4364: color_o = 12'b100000000000;
		13'd4365: color_o = 12'b100000000000;
		13'd4366: color_o = 12'b000000000000;
		13'd4367: color_o = 12'b000000000000;
		13'd4368: color_o = 12'b010000000000;
		13'd4369: color_o = 12'b000000000000;
		13'd4370: color_o = 12'b100000000000;
		13'd4371: color_o = 12'b100000000000;
		13'd4372: color_o = 12'b100000000000;
		13'd4373: color_o = 12'b000000000000;
		13'd4374: color_o = 12'b100000000000;
		13'd4375: color_o = 12'b100000000000;
		13'd4376: color_o = 12'b000000000000;
		13'd4377: color_o = 12'b100000000000;
		13'd4378: color_o = 12'b000000000000;
		13'd4379: color_o = 12'b010000000000;
		13'd4380: color_o = 12'b000000000000;
		13'd4381: color_o = 12'b000000000000;
		13'd4382: color_o = 12'b010001000100;
		13'd4383: color_o = 12'b010001000100;
		13'd4384: color_o = 12'b010001000100;
		13'd4385: color_o = 12'b001101000110;
		13'd4386: color_o = 12'b011110011011;
		13'd4387: color_o = 12'b011110011011;
		13'd4388: color_o = 12'b011101110111;
		13'd4389: color_o = 12'b011101110111;
		13'd4390: color_o = 12'b011110011011;
		13'd4391: color_o = 12'b000000000000;
		13'd4392: color_o = 12'b000000000000;
		13'd4393: color_o = 12'b100000000001;
		13'd4394: color_o = 12'b000000000000;
		13'd4395: color_o = 12'b100000000001;
		13'd4396: color_o = 12'b100000000001;
		13'd4397: color_o = 12'b000000000000;
		13'd4398: color_o = 12'b011101110111;
		13'd4399: color_o = 12'b000011110000;
		13'd4400: color_o = 12'b000011110000;
		13'd4401: color_o = 12'b000011110000;
		13'd4402: color_o = 12'b000011110000;
		13'd4403: color_o = 12'b000011110000;
		13'd4404: color_o = 12'b000011110000;
		13'd4405: color_o = 12'b000011110000;
		13'd4406: color_o = 12'b000011110000;
		13'd4407: color_o = 12'b000011110000;
		13'd4408: color_o = 12'b000011110000;
		13'd4409: color_o = 12'b000011110000;
		13'd4410: color_o = 12'b000011110000;
		13'd4411: color_o = 12'b000011110000;
		13'd4412: color_o = 12'b000011110000;
		13'd4413: color_o = 12'b000011110000;
		13'd4414: color_o = 12'b000011110000;
		13'd4415: color_o = 12'b000011110000;
		13'd4416: color_o = 12'b000011110000;
		13'd4417: color_o = 12'b000011110000;
		13'd4418: color_o = 12'b000011110000;
		13'd4419: color_o = 12'b000000000000;
		13'd4420: color_o = 12'b100000000001;
		13'd4421: color_o = 12'b100000000001;
		13'd4422: color_o = 12'b000000000000;
		13'd4423: color_o = 12'b100000000000;
		13'd4424: color_o = 12'b100000000000;
		13'd4425: color_o = 12'b100000000000;
		13'd4426: color_o = 12'b000000000000;
		13'd4427: color_o = 12'b100000000000;
		13'd4428: color_o = 12'b000000000000;
		13'd4429: color_o = 12'b000000000000;
		13'd4430: color_o = 12'b000000000000;
		13'd4431: color_o = 12'b000000000000;
		13'd4432: color_o = 12'b000000000000;
		13'd4433: color_o = 12'b000000000000;
		13'd4434: color_o = 12'b100000000000;
		13'd4435: color_o = 12'b100000000000;
		13'd4436: color_o = 12'b000000000000;
		13'd4437: color_o = 12'b100000000001;
		13'd4438: color_o = 12'b100000000000;
		13'd4439: color_o = 12'b100000000000;
		13'd4440: color_o = 12'b100000000000;
		13'd4441: color_o = 12'b000000000000;
		13'd4442: color_o = 12'b000000000000;
		13'd4443: color_o = 12'b000000000000;
		13'd4444: color_o = 12'b000000000000;
		13'd4445: color_o = 12'b000000000000;
		13'd4446: color_o = 12'b000000000000;
		13'd4447: color_o = 12'b000000000000;
		13'd4448: color_o = 12'b000000000000;
		13'd4449: color_o = 12'b000000000000;
		13'd4450: color_o = 12'b000000000000;
		13'd4451: color_o = 12'b011101110111;
		13'd4452: color_o = 12'b000000000000;
		13'd4453: color_o = 12'b000000000000;
		13'd4454: color_o = 12'b000000000000;
		13'd4455: color_o = 12'b000000000000;
		13'd4456: color_o = 12'b100000000001;
		13'd4457: color_o = 12'b100000000001;
		13'd4458: color_o = 12'b000000000000;
		13'd4459: color_o = 12'b100000000001;
		13'd4460: color_o = 12'b100000000001;
		13'd4461: color_o = 12'b000000000000;
		13'd4462: color_o = 12'b000000000000;
		13'd4463: color_o = 12'b000011110000;
		13'd4464: color_o = 12'b000011110000;
		13'd4465: color_o = 12'b000011110000;
		13'd4466: color_o = 12'b000011110000;
		13'd4467: color_o = 12'b000011110000;
		13'd4468: color_o = 12'b000011110000;
		13'd4469: color_o = 12'b000011110000;
		13'd4470: color_o = 12'b000011110000;
		13'd4471: color_o = 12'b000011110000;
		13'd4472: color_o = 12'b000011110000;
		13'd4473: color_o = 12'b000011110000;
		13'd4474: color_o = 12'b000011110000;
		13'd4475: color_o = 12'b000011110000;
		13'd4476: color_o = 12'b000011110000;
		13'd4477: color_o = 12'b000011110000;
		13'd4478: color_o = 12'b000011110000;
		13'd4479: color_o = 12'b000011110000;
		13'd4480: color_o = 12'b000011110000;
		13'd4481: color_o = 12'b000011110000;
		13'd4482: color_o = 12'b000000000000;
		13'd4483: color_o = 12'b000000000000;
		13'd4484: color_o = 12'b100000000001;
		13'd4485: color_o = 12'b100000000001;
		13'd4486: color_o = 12'b000000000000;
		13'd4487: color_o = 12'b100000000000;
		13'd4488: color_o = 12'b100000000000;
		13'd4489: color_o = 12'b100000000000;
		13'd4490: color_o = 12'b000000000000;
		13'd4491: color_o = 12'b000000000000;
		13'd4492: color_o = 12'b100000000000;
		13'd4493: color_o = 12'b100000000000;
		13'd4494: color_o = 12'b000000000000;
		13'd4495: color_o = 12'b000000000000;
		13'd4496: color_o = 12'b000000000000;
		13'd4497: color_o = 12'b000000000000;
		13'd4498: color_o = 12'b100000000000;
		13'd4499: color_o = 12'b000000000000;
		13'd4500: color_o = 12'b100000000001;
		13'd4501: color_o = 12'b100000000000;
		13'd4502: color_o = 12'b100000000000;
		13'd4503: color_o = 12'b100000000000;
		13'd4504: color_o = 12'b100000000000;
		13'd4505: color_o = 12'b000000000000;
		13'd4506: color_o = 12'b100000000000;
		13'd4507: color_o = 12'b100000000000;
		13'd4508: color_o = 12'b100000000000;
		13'd4509: color_o = 12'b100000000000;
		13'd4510: color_o = 12'b100000000000;
		13'd4511: color_o = 12'b000000000000;
		13'd4512: color_o = 12'b100000000000;
		13'd4513: color_o = 12'b100000000000;
		13'd4514: color_o = 12'b100000000001;
		13'd4515: color_o = 12'b000000000000;
		13'd4516: color_o = 12'b000000000000;
		13'd4517: color_o = 12'b011101110111;
		13'd4518: color_o = 12'b011101110111;
		13'd4519: color_o = 12'b000000000000;
		13'd4520: color_o = 12'b100000000001;
		13'd4521: color_o = 12'b011101110111;
		13'd4522: color_o = 12'b000000000000;
		13'd4523: color_o = 12'b100000000001;
		13'd4524: color_o = 12'b000000000000;
		13'd4525: color_o = 12'b000011110000;
		13'd4526: color_o = 12'b000011110000;
		13'd4527: color_o = 12'b000011110000;
		13'd4528: color_o = 12'b000011110000;
		13'd4529: color_o = 12'b000011110000;
		13'd4530: color_o = 12'b000011110000;
		13'd4531: color_o = 12'b000011110000;
		13'd4532: color_o = 12'b000011110000;
		13'd4533: color_o = 12'b000011110000;
		13'd4534: color_o = 12'b000011110000;
		13'd4535: color_o = 12'b000011110000;
		13'd4536: color_o = 12'b000011110000;
		13'd4537: color_o = 12'b000011110000;
		13'd4538: color_o = 12'b000011110000;
		13'd4539: color_o = 12'b000011110000;
		13'd4540: color_o = 12'b000011110000;
		13'd4541: color_o = 12'b000011110000;
		13'd4542: color_o = 12'b000011110000;
		13'd4543: color_o = 12'b000011110000;
		13'd4544: color_o = 12'b000011110000;
		13'd4545: color_o = 12'b000011110000;
		13'd4546: color_o = 12'b000000000000;
		13'd4547: color_o = 12'b000000000000;
		13'd4548: color_o = 12'b100000000001;
		13'd4549: color_o = 12'b100000000001;
		13'd4550: color_o = 12'b000000000000;
		13'd4551: color_o = 12'b100000000000;
		13'd4552: color_o = 12'b100000000000;
		13'd4553: color_o = 12'b100000000000;
		13'd4554: color_o = 12'b100000000000;
		13'd4555: color_o = 12'b100000000000;
		13'd4556: color_o = 12'b000000000000;
		13'd4557: color_o = 12'b100000000000;
		13'd4558: color_o = 12'b100000000000;
		13'd4559: color_o = 12'b100000000000;
		13'd4560: color_o = 12'b100000000000;
		13'd4561: color_o = 12'b100000000000;
		13'd4562: color_o = 12'b100000000000;
		13'd4563: color_o = 12'b100000000000;
		13'd4564: color_o = 12'b100000000000;
		13'd4565: color_o = 12'b100000000000;
		13'd4566: color_o = 12'b100000000000;
		13'd4567: color_o = 12'b100000000000;
		13'd4568: color_o = 12'b100000000000;
		13'd4569: color_o = 12'b100000000000;
		13'd4570: color_o = 12'b100000000000;
		13'd4571: color_o = 12'b100000000000;
		13'd4572: color_o = 12'b100000000000;
		13'd4573: color_o = 12'b100000000000;
		13'd4574: color_o = 12'b100000000000;
		13'd4575: color_o = 12'b100000000000;
		13'd4576: color_o = 12'b100000000000;
		13'd4577: color_o = 12'b100000000000;
		13'd4578: color_o = 12'b100000000001;
		13'd4579: color_o = 12'b000000000000;
		13'd4580: color_o = 12'b000000000000;
		13'd4581: color_o = 12'b011101110111;
		13'd4582: color_o = 12'b011101110111;
		13'd4583: color_o = 12'b011101110111;
		13'd4584: color_o = 12'b011101110111;
		13'd4585: color_o = 12'b011101110111;
		13'd4586: color_o = 12'b000000000000;
		13'd4587: color_o = 12'b000000000000;
		13'd4588: color_o = 12'b000011110000;
		13'd4589: color_o = 12'b000011110000;
		13'd4590: color_o = 12'b000011110000;
		13'd4591: color_o = 12'b000011110000;
		13'd4592: color_o = 12'b000011110000;
		13'd4593: color_o = 12'b000011110000;
		13'd4594: color_o = 12'b000011110000;
		13'd4595: color_o = 12'b000011110000;
		13'd4596: color_o = 12'b000011110000;
		13'd4597: color_o = 12'b000011110000;
		13'd4598: color_o = 12'b000011110000;
		13'd4599: color_o = 12'b000011110000;
		13'd4600: color_o = 12'b000011110000;
		13'd4601: color_o = 12'b000011110000;
		13'd4602: color_o = 12'b000011110000;
		13'd4603: color_o = 12'b000011110000;
		13'd4604: color_o = 12'b000011110000;
		13'd4605: color_o = 12'b000011110000;
		13'd4606: color_o = 12'b000011110000;
		13'd4607: color_o = 12'b000011110000;
		13'd4608: color_o = 12'b000011110000;
		13'd4609: color_o = 12'b000011110000;
		13'd4610: color_o = 12'b000000000000;
		13'd4611: color_o = 12'b000000000000;
		13'd4612: color_o = 12'b100000000001;
		13'd4613: color_o = 12'b100000000001;
		13'd4614: color_o = 12'b000000000000;
		13'd4615: color_o = 12'b000000000000;
		13'd4616: color_o = 12'b100000000000;
		13'd4617: color_o = 12'b100000000000;
		13'd4618: color_o = 12'b100000000000;
		13'd4619: color_o = 12'b100000000000;
		13'd4620: color_o = 12'b000000000000;
		13'd4621: color_o = 12'b000000000000;
		13'd4622: color_o = 12'b000000000000;
		13'd4623: color_o = 12'b000000000000;
		13'd4624: color_o = 12'b100000000000;
		13'd4625: color_o = 12'b000000000000;
		13'd4626: color_o = 12'b100000000000;
		13'd4627: color_o = 12'b100000000000;
		13'd4628: color_o = 12'b100000000000;
		13'd4629: color_o = 12'b100000000000;
		13'd4630: color_o = 12'b100000000000;
		13'd4631: color_o = 12'b100000000000;
		13'd4632: color_o = 12'b100000000000;
		13'd4633: color_o = 12'b000000000000;
		13'd4634: color_o = 12'b000000000000;
		13'd4635: color_o = 12'b100000000000;
		13'd4636: color_o = 12'b100000000000;
		13'd4637: color_o = 12'b100000000000;
		13'd4638: color_o = 12'b100000000000;
		13'd4639: color_o = 12'b000000000000;
		13'd4640: color_o = 12'b000000000000;
		13'd4641: color_o = 12'b100000000000;
		13'd4642: color_o = 12'b100000000001;
		13'd4643: color_o = 12'b000000000000;
		13'd4644: color_o = 12'b100000000001;
		13'd4645: color_o = 12'b000000000000;
		13'd4646: color_o = 12'b000000000000;
		13'd4647: color_o = 12'b011101110111;
		13'd4648: color_o = 12'b011101110111;
		13'd4649: color_o = 12'b011101110111;
		13'd4650: color_o = 12'b000000000000;
		13'd4651: color_o = 12'b000000000000;
		13'd4652: color_o = 12'b000011110000;
		13'd4653: color_o = 12'b000011110000;
		13'd4654: color_o = 12'b000011110000;
		13'd4655: color_o = 12'b000011110000;
		13'd4656: color_o = 12'b000011110000;
		13'd4657: color_o = 12'b000011110000;
		13'd4658: color_o = 12'b000011110000;
		13'd4659: color_o = 12'b000011110000;
		13'd4660: color_o = 12'b000011110000;
		13'd4661: color_o = 12'b000011110000;
		13'd4662: color_o = 12'b000011110000;
		13'd4663: color_o = 12'b000011110000;
		13'd4664: color_o = 12'b000011110000;
		13'd4665: color_o = 12'b000011110000;
		13'd4666: color_o = 12'b000011110000;
		13'd4667: color_o = 12'b000011110000;
		13'd4668: color_o = 12'b000011110000;
		13'd4669: color_o = 12'b000011110000;
		13'd4670: color_o = 12'b000011110000;
		13'd4671: color_o = 12'b000011110000;
		13'd4672: color_o = 12'b000011110000;
		13'd4673: color_o = 12'b000011110000;
		13'd4674: color_o = 12'b000000000000;
		13'd4675: color_o = 12'b000000000000;
		13'd4676: color_o = 12'b100000000001;
		13'd4677: color_o = 12'b100000000001;
		13'd4678: color_o = 12'b100000000001;
		13'd4679: color_o = 12'b000000000000;
		13'd4680: color_o = 12'b100000000000;
		13'd4681: color_o = 12'b000000000000;
		13'd4682: color_o = 12'b100000000000;
		13'd4683: color_o = 12'b000000000000;
		13'd4684: color_o = 12'b100000000000;
		13'd4685: color_o = 12'b010000000000;
		13'd4686: color_o = 12'b010000000000;
		13'd4687: color_o = 12'b000000000000;
		13'd4688: color_o = 12'b010000000000;
		13'd4689: color_o = 12'b100000000000;
		13'd4690: color_o = 12'b010000000000;
		13'd4691: color_o = 12'b100000000000;
		13'd4692: color_o = 12'b100000000000;
		13'd4693: color_o = 12'b100000000000;
		13'd4694: color_o = 12'b100000000000;
		13'd4695: color_o = 12'b100000000000;
		13'd4696: color_o = 12'b000000000000;
		13'd4697: color_o = 12'b100000000000;
		13'd4698: color_o = 12'b100000000000;
		13'd4699: color_o = 12'b000000000000;
		13'd4700: color_o = 12'b100000000000;
		13'd4701: color_o = 12'b000000000000;
		13'd4702: color_o = 12'b000000000000;
		13'd4703: color_o = 12'b100000000000;
		13'd4704: color_o = 12'b100000000000;
		13'd4705: color_o = 12'b100000000000;
		13'd4706: color_o = 12'b100000000000;
		13'd4707: color_o = 12'b010000000000;
		13'd4708: color_o = 12'b000000000000;
		13'd4709: color_o = 12'b000011110000;
		13'd4710: color_o = 12'b000000000000;
		13'd4711: color_o = 12'b000000000000;
		13'd4712: color_o = 12'b011101110111;
		13'd4713: color_o = 12'b000000000000;
		13'd4714: color_o = 12'b000000000000;
		13'd4715: color_o = 12'b000011110000;
		13'd4716: color_o = 12'b000011110000;
		13'd4717: color_o = 12'b000011110000;
		13'd4718: color_o = 12'b000011110000;
		13'd4719: color_o = 12'b000011110000;
		13'd4720: color_o = 12'b000011110000;
		13'd4721: color_o = 12'b000011110000;
		13'd4722: color_o = 12'b000011110000;
		13'd4723: color_o = 12'b000011110000;
		13'd4724: color_o = 12'b000011110000;
		13'd4725: color_o = 12'b000011110000;
		13'd4726: color_o = 12'b000011110000;
		13'd4727: color_o = 12'b000011110000;
		13'd4728: color_o = 12'b000011110000;
		13'd4729: color_o = 12'b000011110000;
		13'd4730: color_o = 12'b000011110000;
		13'd4731: color_o = 12'b000011110000;
		13'd4732: color_o = 12'b000011110000;
		13'd4733: color_o = 12'b000011110000;
		13'd4734: color_o = 12'b000011110000;
		13'd4735: color_o = 12'b000011110000;
		13'd4736: color_o = 12'b000011110000;
		13'd4737: color_o = 12'b000000000000;
		13'd4738: color_o = 12'b000000000000;
		13'd4739: color_o = 12'b010000000000;
		13'd4740: color_o = 12'b100000000001;
		13'd4741: color_o = 12'b100000000001;
		13'd4742: color_o = 12'b100000000001;
		13'd4743: color_o = 12'b000000000000;
		13'd4744: color_o = 12'b100000000000;
		13'd4745: color_o = 12'b100000000000;
		13'd4746: color_o = 12'b100000000000;
		13'd4747: color_o = 12'b100000000000;
		13'd4748: color_o = 12'b100000000000;
		13'd4749: color_o = 12'b100000000000;
		13'd4750: color_o = 12'b010000000000;
		13'd4751: color_o = 12'b000000000000;
		13'd4752: color_o = 12'b000000000000;
		13'd4753: color_o = 12'b010000000000;
		13'd4754: color_o = 12'b100000000001;
		13'd4755: color_o = 12'b010000000000;
		13'd4756: color_o = 12'b100000000000;
		13'd4757: color_o = 12'b100000000000;
		13'd4758: color_o = 12'b100000000000;
		13'd4759: color_o = 12'b100000000000;
		13'd4760: color_o = 12'b100000000000;
		13'd4761: color_o = 12'b100000000000;
		13'd4762: color_o = 12'b100000000000;
		13'd4763: color_o = 12'b100000000000;
		13'd4764: color_o = 12'b000000000000;
		13'd4765: color_o = 12'b100000000000;
		13'd4766: color_o = 12'b100000000000;
		13'd4767: color_o = 12'b100000000000;
		13'd4768: color_o = 12'b010000000000;
		13'd4769: color_o = 12'b010000000000;
		13'd4770: color_o = 12'b000000000000;
		13'd4771: color_o = 12'b000000000000;
		13'd4772: color_o = 12'b000011110000;
		13'd4773: color_o = 12'b000011110000;
		13'd4774: color_o = 12'b000011110000;
		13'd4775: color_o = 12'b000000000000;
		13'd4776: color_o = 12'b011101110111;
		13'd4777: color_o = 12'b000011110000;
		13'd4778: color_o = 12'b000011110000;
		13'd4779: color_o = 12'b000011110000;
		13'd4780: color_o = 12'b000011110000;
		13'd4781: color_o = 12'b000011110000;
		13'd4782: color_o = 12'b000011110000;
		13'd4783: color_o = 12'b000011110000;
		13'd4784: color_o = 12'b000011110000;
		13'd4785: color_o = 12'b000011110000;
		13'd4786: color_o = 12'b000011110000;
		13'd4787: color_o = 12'b000011110000;
		13'd4788: color_o = 12'b000011110000;
		13'd4789: color_o = 12'b000011110000;
		13'd4790: color_o = 12'b000011110000;
		13'd4791: color_o = 12'b000011110000;
		13'd4792: color_o = 12'b000011110000;
		13'd4793: color_o = 12'b000011110000;
		13'd4794: color_o = 12'b000011110000;
		13'd4795: color_o = 12'b000011110000;
		13'd4796: color_o = 12'b000011110000;
		13'd4797: color_o = 12'b000011110000;
		13'd4798: color_o = 12'b000011110000;
		13'd4799: color_o = 12'b000011110000;
		13'd4800: color_o = 12'b000011110000;
		13'd4801: color_o = 12'b000000000000;
		13'd4802: color_o = 12'b000000000000;
		13'd4803: color_o = 12'b010000000000;
		13'd4804: color_o = 12'b100000000001;
		13'd4805: color_o = 12'b100000000001;
		13'd4806: color_o = 12'b100000000001;
		13'd4807: color_o = 12'b000000000000;
		13'd4808: color_o = 12'b100000000000;
		13'd4809: color_o = 12'b000000000000;
		13'd4810: color_o = 12'b100000000000;
		13'd4811: color_o = 12'b100000000000;
		13'd4812: color_o = 12'b100000000001;
		13'd4813: color_o = 12'b100000000000;
		13'd4814: color_o = 12'b010000000000;
		13'd4815: color_o = 12'b010000000000;
		13'd4816: color_o = 12'b000000000000;
		13'd4817: color_o = 12'b000000000000;
		13'd4818: color_o = 12'b010000000000;
		13'd4819: color_o = 12'b100000000000;
		13'd4820: color_o = 12'b010000000000;
		13'd4821: color_o = 12'b100000000001;
		13'd4822: color_o = 12'b100000000001;
		13'd4823: color_o = 12'b000000000000;
		13'd4824: color_o = 12'b100000000000;
		13'd4825: color_o = 12'b100000000000;
		13'd4826: color_o = 12'b100000000000;
		13'd4827: color_o = 12'b100000000000;
		13'd4828: color_o = 12'b000000000000;
		13'd4829: color_o = 12'b010000000000;
		13'd4830: color_o = 12'b010000000000;
		13'd4831: color_o = 12'b010000000000;
		13'd4832: color_o = 12'b000000000000;
		13'd4833: color_o = 12'b000000000000;
		13'd4834: color_o = 12'b000011110000;
		13'd4835: color_o = 12'b000011110000;
		13'd4836: color_o = 12'b000011110000;
		13'd4837: color_o = 12'b000011110000;
		13'd4838: color_o = 12'b000011110000;
		13'd4839: color_o = 12'b000000000000;
		13'd4840: color_o = 12'b000000000000;
		13'd4841: color_o = 12'b000011110000;
		13'd4842: color_o = 12'b000011110000;
		13'd4843: color_o = 12'b000011110000;
		13'd4844: color_o = 12'b000011110000;
		13'd4845: color_o = 12'b000011110000;
		13'd4846: color_o = 12'b000011110000;
		13'd4847: color_o = 12'b000011110000;
		13'd4848: color_o = 12'b000011110000;
		13'd4849: color_o = 12'b000011110000;
		13'd4850: color_o = 12'b000011110000;
		13'd4851: color_o = 12'b000011110000;
		13'd4852: color_o = 12'b000011110000;
		13'd4853: color_o = 12'b000011110000;
		13'd4854: color_o = 12'b000011110000;
		13'd4855: color_o = 12'b000011110000;
		13'd4856: color_o = 12'b000011110000;
		13'd4857: color_o = 12'b000011110000;
		13'd4858: color_o = 12'b000011110000;
		13'd4859: color_o = 12'b000011110000;
		13'd4860: color_o = 12'b000011110000;
		13'd4861: color_o = 12'b000011110000;
		13'd4862: color_o = 12'b000011110000;
		13'd4863: color_o = 12'b000011110000;
		13'd4864: color_o = 12'b000011110000;
		13'd4865: color_o = 12'b000000000000;
		13'd4866: color_o = 12'b000000000000;
		13'd4867: color_o = 12'b010000000000;
		13'd4868: color_o = 12'b100000000001;
		13'd4869: color_o = 12'b100000000001;
		13'd4870: color_o = 12'b100000000001;
		13'd4871: color_o = 12'b000000000000;
		13'd4872: color_o = 12'b000000000000;
		13'd4873: color_o = 12'b000000000000;
		13'd4874: color_o = 12'b100000000001;
		13'd4875: color_o = 12'b100000000001;
		13'd4876: color_o = 12'b100000000001;
		13'd4877: color_o = 12'b100000000000;
		13'd4878: color_o = 12'b100000000000;
		13'd4879: color_o = 12'b010000000000;
		13'd4880: color_o = 12'b010000000000;
		13'd4881: color_o = 12'b000000000000;
		13'd4882: color_o = 12'b000000000000;
		13'd4883: color_o = 12'b010000000000;
		13'd4884: color_o = 12'b010000000000;
		13'd4885: color_o = 12'b010000000000;
		13'd4886: color_o = 12'b010000000000;
		13'd4887: color_o = 12'b010000000000;
		13'd4888: color_o = 12'b000000000000;
		13'd4889: color_o = 12'b100000000000;
		13'd4890: color_o = 12'b100000000000;
		13'd4891: color_o = 12'b010000000000;
		13'd4892: color_o = 12'b000000000000;
		13'd4893: color_o = 12'b000000000000;
		13'd4894: color_o = 12'b000000000000;
		13'd4895: color_o = 12'b000000000000;
		13'd4896: color_o = 12'b000011110000;
		13'd4897: color_o = 12'b000011110000;
		13'd4898: color_o = 12'b000011110000;
		13'd4899: color_o = 12'b000011110000;
		13'd4900: color_o = 12'b000011110000;
		13'd4901: color_o = 12'b000011110000;
		13'd4902: color_o = 12'b000011110000;
		13'd4903: color_o = 12'b000011110000;
		13'd4904: color_o = 12'b000000000000;
		13'd4905: color_o = 12'b000011110000;
		13'd4906: color_o = 12'b000011110000;
		13'd4907: color_o = 12'b000011110000;
		13'd4908: color_o = 12'b000011110000;
		13'd4909: color_o = 12'b000011110000;
		13'd4910: color_o = 12'b000011110000;
		13'd4911: color_o = 12'b000011110000;
		13'd4912: color_o = 12'b000011110000;
		13'd4913: color_o = 12'b000011110000;
		13'd4914: color_o = 12'b000011110000;
		13'd4915: color_o = 12'b000011110000;
		13'd4916: color_o = 12'b000011110000;
		13'd4917: color_o = 12'b000011110000;
		13'd4918: color_o = 12'b000011110000;
		13'd4919: color_o = 12'b000011110000;
		13'd4920: color_o = 12'b000011110000;
		13'd4921: color_o = 12'b000011110000;
		13'd4922: color_o = 12'b000011110000;
		13'd4923: color_o = 12'b000011110000;
		13'd4924: color_o = 12'b000011110000;
		13'd4925: color_o = 12'b000011110000;
		13'd4926: color_o = 12'b000011110000;
		13'd4927: color_o = 12'b000011110000;
		13'd4928: color_o = 12'b000011110000;
		13'd4929: color_o = 12'b000000000000;
		13'd4930: color_o = 12'b000000000000;
		13'd4931: color_o = 12'b010000000000;
		13'd4932: color_o = 12'b100000000001;
		13'd4933: color_o = 12'b100000000001;
		13'd4934: color_o = 12'b100000000001;
		13'd4935: color_o = 12'b000000000000;
		13'd4936: color_o = 12'b000000000000;
		13'd4937: color_o = 12'b100000000001;
		13'd4938: color_o = 12'b100000000001;
		13'd4939: color_o = 12'b100000000001;
		13'd4940: color_o = 12'b100000000001;
		13'd4941: color_o = 12'b100000000001;
		13'd4942: color_o = 12'b100000000000;
		13'd4943: color_o = 12'b100000000000;
		13'd4944: color_o = 12'b100000000000;
		13'd4945: color_o = 12'b100000000000;
		13'd4946: color_o = 12'b000000000000;
		13'd4947: color_o = 12'b000000000000;
		13'd4948: color_o = 12'b000000000000;
		13'd4949: color_o = 12'b000000000000;
		13'd4950: color_o = 12'b000000000000;
		13'd4951: color_o = 12'b000000000000;
		13'd4952: color_o = 12'b000000000000;
		13'd4953: color_o = 12'b010000000000;
		13'd4954: color_o = 12'b010000000000;
		13'd4955: color_o = 12'b000000000000;
		13'd4956: color_o = 12'b000000000000;
		13'd4957: color_o = 12'b000000000000;
		13'd4958: color_o = 12'b000011110000;
		13'd4959: color_o = 12'b000011110000;
		13'd4960: color_o = 12'b000011110000;
		13'd4961: color_o = 12'b000011110000;
		13'd4962: color_o = 12'b000011110000;
		13'd4963: color_o = 12'b000011110000;
		13'd4964: color_o = 12'b000011110000;
		13'd4965: color_o = 12'b000011110000;
		13'd4966: color_o = 12'b000011110000;
		13'd4967: color_o = 12'b000011110000;
		13'd4968: color_o = 12'b000011110000;
		13'd4969: color_o = 12'b000011110000;
		13'd4970: color_o = 12'b000011110000;
		13'd4971: color_o = 12'b000011110000;
		13'd4972: color_o = 12'b000011110000;
		13'd4973: color_o = 12'b000011110000;
		13'd4974: color_o = 12'b000011110000;
		13'd4975: color_o = 12'b000011110000;
		13'd4976: color_o = 12'b000011110000;
		13'd4977: color_o = 12'b000011110000;
		13'd4978: color_o = 12'b000011110000;
		13'd4979: color_o = 12'b000011110000;
		13'd4980: color_o = 12'b000011110000;
		13'd4981: color_o = 12'b000011110000;
		13'd4982: color_o = 12'b000011110000;
		13'd4983: color_o = 12'b000011110000;
		13'd4984: color_o = 12'b000011110000;
		13'd4985: color_o = 12'b000011110000;
		13'd4986: color_o = 12'b000011110000;
		13'd4987: color_o = 12'b000011110000;
		13'd4988: color_o = 12'b000011110000;
		13'd4989: color_o = 12'b000011110000;
		13'd4990: color_o = 12'b000011110000;
		13'd4991: color_o = 12'b000011110000;
		13'd4992: color_o = 12'b000011110000;
		13'd4993: color_o = 12'b000000000000;
		13'd4994: color_o = 12'b000000000000;
		13'd4995: color_o = 12'b010000000000;
		13'd4996: color_o = 12'b010000000000;
		13'd4997: color_o = 12'b100000000001;
		13'd4998: color_o = 12'b000000000000;
		13'd4999: color_o = 12'b000000000000;
		13'd5000: color_o = 12'b000000000000;
		13'd5001: color_o = 12'b000000000000;
		13'd5002: color_o = 12'b000000000000;
		13'd5003: color_o = 12'b100000000001;
		13'd5004: color_o = 12'b100000000001;
		13'd5005: color_o = 12'b010000000000;
		13'd5006: color_o = 12'b010000000000;
		13'd5007: color_o = 12'b010000000000;
		13'd5008: color_o = 12'b010000000000;
		13'd5009: color_o = 12'b100000000000;
		13'd5010: color_o = 12'b100000000000;
		13'd5011: color_o = 12'b010000000000;
		13'd5012: color_o = 12'b010000000000;
		13'd5013: color_o = 12'b010000000000;
		13'd5014: color_o = 12'b010000000000;
		13'd5015: color_o = 12'b010000000000;
		13'd5016: color_o = 12'b010000000000;
		13'd5017: color_o = 12'b000000000000;
		13'd5018: color_o = 12'b000000000000;
		13'd5019: color_o = 12'b100000000001;
		13'd5020: color_o = 12'b000000000000;
		13'd5021: color_o = 12'b000011110000;
		13'd5022: color_o = 12'b000011110000;
		13'd5023: color_o = 12'b000011110000;
		13'd5024: color_o = 12'b000011110000;
		13'd5025: color_o = 12'b000011110000;
		13'd5026: color_o = 12'b000011110000;
		13'd5027: color_o = 12'b000011110000;
		13'd5028: color_o = 12'b000011110000;
		13'd5029: color_o = 12'b000011110000;
		13'd5030: color_o = 12'b000011110000;
		13'd5031: color_o = 12'b000011110000;
		13'd5032: color_o = 12'b000011110000;
		13'd5033: color_o = 12'b000011110000;
		13'd5034: color_o = 12'b000011110000;
		13'd5035: color_o = 12'b000011110000;
		13'd5036: color_o = 12'b000011110000;
		13'd5037: color_o = 12'b000011110000;
		13'd5038: color_o = 12'b000011110000;
		13'd5039: color_o = 12'b000011110000;
		13'd5040: color_o = 12'b000011110000;
		13'd5041: color_o = 12'b000011110000;
		13'd5042: color_o = 12'b000011110000;
		13'd5043: color_o = 12'b000011110000;
		13'd5044: color_o = 12'b000011110000;
		13'd5045: color_o = 12'b000011110000;
		13'd5046: color_o = 12'b000011110000;
		13'd5047: color_o = 12'b000011110000;
		13'd5048: color_o = 12'b000011110000;
		13'd5049: color_o = 12'b000011110000;
		13'd5050: color_o = 12'b000011110000;
		13'd5051: color_o = 12'b000011110000;
		13'd5052: color_o = 12'b000011110000;
		13'd5053: color_o = 12'b000011110000;
		13'd5054: color_o = 12'b000011110000;
		13'd5055: color_o = 12'b000011110000;
		13'd5056: color_o = 12'b000011110000;
		13'd5057: color_o = 12'b000000000000;
		13'd5058: color_o = 12'b000000000000;
		13'd5059: color_o = 12'b010000000000;
		13'd5060: color_o = 12'b010000000000;
		13'd5061: color_o = 12'b000000000000;
		13'd5062: color_o = 12'b000000000000;
		13'd5063: color_o = 12'b100000000000;
		13'd5064: color_o = 12'b000000000000;
		13'd5065: color_o = 12'b000000000000;
		13'd5066: color_o = 12'b000000000000;
		13'd5067: color_o = 12'b100000000001;
		13'd5068: color_o = 12'b100000000001;
		13'd5069: color_o = 12'b100000000001;
		13'd5070: color_o = 12'b100000000001;
		13'd5071: color_o = 12'b100000000001;
		13'd5072: color_o = 12'b010000000000;
		13'd5073: color_o = 12'b010000000000;
		13'd5074: color_o = 12'b010000000000;
		13'd5075: color_o = 12'b010000000000;
		13'd5076: color_o = 12'b010000000000;
		13'd5077: color_o = 12'b100000000001;
		13'd5078: color_o = 12'b100000000001;
		13'd5079: color_o = 12'b100000000000;
		13'd5080: color_o = 12'b100000000000;
		13'd5081: color_o = 12'b100000000000;
		13'd5082: color_o = 12'b100000000000;
		13'd5083: color_o = 12'b100000000000;
		13'd5084: color_o = 12'b000000000000;
		13'd5085: color_o = 12'b000011110000;
		13'd5086: color_o = 12'b000011110000;
		13'd5087: color_o = 12'b000011110000;
		13'd5088: color_o = 12'b000011110000;
		13'd5089: color_o = 12'b000011110000;
		13'd5090: color_o = 12'b000011110000;
		13'd5091: color_o = 12'b000011110000;
		13'd5092: color_o = 12'b000011110000;
		13'd5093: color_o = 12'b000011110000;
		13'd5094: color_o = 12'b000011110000;
		13'd5095: color_o = 12'b000011110000;
		13'd5096: color_o = 12'b000011110000;
		13'd5097: color_o = 12'b000011110000;
		13'd5098: color_o = 12'b000011110000;
		13'd5099: color_o = 12'b000011110000;
		13'd5100: color_o = 12'b000011110000;
		13'd5101: color_o = 12'b000011110000;
		13'd5102: color_o = 12'b000011110000;
		13'd5103: color_o = 12'b000011110000;
		13'd5104: color_o = 12'b000011110000;
		13'd5105: color_o = 12'b000011110000;
		13'd5106: color_o = 12'b000011110000;
		13'd5107: color_o = 12'b000011110000;
		13'd5108: color_o = 12'b000011110000;
		13'd5109: color_o = 12'b000011110000;
		13'd5110: color_o = 12'b000011110000;
		13'd5111: color_o = 12'b000011110000;
		13'd5112: color_o = 12'b000011110000;
		13'd5113: color_o = 12'b000011110000;
		13'd5114: color_o = 12'b000011110000;
		13'd5115: color_o = 12'b000011110000;
		13'd5116: color_o = 12'b000011110000;
		13'd5117: color_o = 12'b000011110000;
		13'd5118: color_o = 12'b000011110000;
		13'd5119: color_o = 12'b000011110000;
		13'd5120: color_o = 12'b000011110000;
		13'd5121: color_o = 12'b000000000000;
		13'd5122: color_o = 12'b000000000000;
		13'd5123: color_o = 12'b010000000000;
		13'd5124: color_o = 12'b000000000000;
		13'd5125: color_o = 12'b000000000000;
		13'd5126: color_o = 12'b100000000000;
		13'd5127: color_o = 12'b100000000000;
		13'd5128: color_o = 12'b000000000000;
		13'd5129: color_o = 12'b000000000000;
		13'd5130: color_o = 12'b000000000000;
		13'd5131: color_o = 12'b000000000000;
		13'd5132: color_o = 12'b100000000001;
		13'd5133: color_o = 12'b100000000001;
		13'd5134: color_o = 12'b100000000001;
		13'd5135: color_o = 12'b100000000001;
		13'd5136: color_o = 12'b100000000000;
		13'd5137: color_o = 12'b100000000001;
		13'd5138: color_o = 12'b100000000001;
		13'd5139: color_o = 12'b100000000001;
		13'd5140: color_o = 12'b100000000000;
		13'd5141: color_o = 12'b100000000001;
		13'd5142: color_o = 12'b100000000000;
		13'd5143: color_o = 12'b100000000000;
		13'd5144: color_o = 12'b100000000000;
		13'd5145: color_o = 12'b000000000000;
		13'd5146: color_o = 12'b000000000000;
		13'd5147: color_o = 12'b000000000000;
		13'd5148: color_o = 12'b000000000000;
		13'd5149: color_o = 12'b000011110000;
		13'd5150: color_o = 12'b000011110000;
		13'd5151: color_o = 12'b000011110000;
		13'd5152: color_o = 12'b000011110000;
		13'd5153: color_o = 12'b000011110000;
		13'd5154: color_o = 12'b000011110000;
		13'd5155: color_o = 12'b000011110000;
		13'd5156: color_o = 12'b000011110000;
		13'd5157: color_o = 12'b000011110000;
		13'd5158: color_o = 12'b000011110000;
		13'd5159: color_o = 12'b000011110000;
		13'd5160: color_o = 12'b000011110000;
		13'd5161: color_o = 12'b000011110000;
		13'd5162: color_o = 12'b000011110000;
		13'd5163: color_o = 12'b000011110000;
		13'd5164: color_o = 12'b000011110000;
		13'd5165: color_o = 12'b000011110000;
		13'd5166: color_o = 12'b000011110000;
		13'd5167: color_o = 12'b000011110000;
		13'd5168: color_o = 12'b000011110000;
		13'd5169: color_o = 12'b000011110000;
		13'd5170: color_o = 12'b000011110000;
		13'd5171: color_o = 12'b000011110000;
		13'd5172: color_o = 12'b000011110000;
		13'd5173: color_o = 12'b000011110000;
		13'd5174: color_o = 12'b000011110000;
		13'd5175: color_o = 12'b000011110000;
		13'd5176: color_o = 12'b000011110000;
		13'd5177: color_o = 12'b000011110000;
		13'd5178: color_o = 12'b000011110000;
		13'd5179: color_o = 12'b000011110000;
		13'd5180: color_o = 12'b000011110000;
		13'd5181: color_o = 12'b000011110000;
		13'd5182: color_o = 12'b000011110000;
		13'd5183: color_o = 12'b000011110000;
		13'd5184: color_o = 12'b000011110000;
		13'd5185: color_o = 12'b000000000000;
		13'd5186: color_o = 12'b000000000000;
		13'd5187: color_o = 12'b000000000000;
		13'd5188: color_o = 12'b000000000000;
		13'd5189: color_o = 12'b000000000000;
		13'd5190: color_o = 12'b100000000001;
		13'd5191: color_o = 12'b100000000001;
		13'd5192: color_o = 12'b000000000000;
		13'd5193: color_o = 12'b000000000000;
		13'd5194: color_o = 12'b100000000000;
		13'd5195: color_o = 12'b000000000000;
		13'd5196: color_o = 12'b000000000000;
		13'd5197: color_o = 12'b000000000000;
		13'd5198: color_o = 12'b000000000000;
		13'd5199: color_o = 12'b100000000000;
		13'd5200: color_o = 12'b100000000001;
		13'd5201: color_o = 12'b100000000001;
		13'd5202: color_o = 12'b100000000001;
		13'd5203: color_o = 12'b100000000001;
		13'd5204: color_o = 12'b100000000001;
		13'd5205: color_o = 12'b100000000000;
		13'd5206: color_o = 12'b100000000000;
		13'd5207: color_o = 12'b100000000000;
		13'd5208: color_o = 12'b000000000000;
		13'd5209: color_o = 12'b000000000000;
		13'd5210: color_o = 12'b100000000000;
		13'd5211: color_o = 12'b100000000000;
		13'd5212: color_o = 12'b000000000000;
		13'd5213: color_o = 12'b000011110000;
		13'd5214: color_o = 12'b000011110000;
		13'd5215: color_o = 12'b000011110000;
		13'd5216: color_o = 12'b000011110000;
		13'd5217: color_o = 12'b000011110000;
		13'd5218: color_o = 12'b000011110000;
		13'd5219: color_o = 12'b000011110000;
		13'd5220: color_o = 12'b000011110000;
		13'd5221: color_o = 12'b000011110000;
		13'd5222: color_o = 12'b000011110000;
		13'd5223: color_o = 12'b000011110000;
		13'd5224: color_o = 12'b000011110000;
		13'd5225: color_o = 12'b000011110000;
		13'd5226: color_o = 12'b000011110000;
		13'd5227: color_o = 12'b000011110000;
		13'd5228: color_o = 12'b000011110000;
		13'd5229: color_o = 12'b000011110000;
		13'd5230: color_o = 12'b000011110000;
		13'd5231: color_o = 12'b000011110000;
		13'd5232: color_o = 12'b000011110000;
		13'd5233: color_o = 12'b000011110000;
		13'd5234: color_o = 12'b000011110000;
		13'd5235: color_o = 12'b000011110000;
		13'd5236: color_o = 12'b000011110000;
		13'd5237: color_o = 12'b000011110000;
		13'd5238: color_o = 12'b000011110000;
		13'd5239: color_o = 12'b000011110000;
		13'd5240: color_o = 12'b000011110000;
		13'd5241: color_o = 12'b000011110000;
		13'd5242: color_o = 12'b000011110000;
		13'd5243: color_o = 12'b000011110000;
		13'd5244: color_o = 12'b000011110000;
		13'd5245: color_o = 12'b000011110000;
		13'd5246: color_o = 12'b000011110000;
		13'd5247: color_o = 12'b000011110000;
		13'd5248: color_o = 12'b000011110000;
		13'd5249: color_o = 12'b000011110000;
		13'd5250: color_o = 12'b000011110000;
		13'd5251: color_o = 12'b000011110000;
		13'd5252: color_o = 12'b000000000000;
		13'd5253: color_o = 12'b000000000000;
		13'd5254: color_o = 12'b000000000000;
		13'd5255: color_o = 12'b000000000000;
		13'd5256: color_o = 12'b000000000000;
		13'd5257: color_o = 12'b000000000000;
		13'd5258: color_o = 12'b000000000000;
		13'd5259: color_o = 12'b000000000000;
		13'd5260: color_o = 12'b100000000000;
		13'd5261: color_o = 12'b000000000000;
		13'd5262: color_o = 12'b000000000000;
		13'd5263: color_o = 12'b000000000000;
		13'd5264: color_o = 12'b000000000000;
		13'd5265: color_o = 12'b000000000000;
		13'd5266: color_o = 12'b000000000000;
		13'd5267: color_o = 12'b000000000000;
		13'd5268: color_o = 12'b100000000001;
		13'd5269: color_o = 12'b100000000001;
		13'd5270: color_o = 12'b000000000000;
		13'd5271: color_o = 12'b000000000000;
		13'd5272: color_o = 12'b000000000000;
		13'd5273: color_o = 12'b000000000000;
		13'd5274: color_o = 12'b000000000000;
		13'd5275: color_o = 12'b000000000000;
		13'd5276: color_o = 12'b000011110000;
		13'd5277: color_o = 12'b000011110000;
		13'd5278: color_o = 12'b000011110000;
		13'd5279: color_o = 12'b000011110000;
		13'd5280: color_o = 12'b000011110000;
		13'd5281: color_o = 12'b000011110000;
		13'd5282: color_o = 12'b000011110000;
		13'd5283: color_o = 12'b000011110000;
		13'd5284: color_o = 12'b000011110000;
		13'd5285: color_o = 12'b000011110000;
		13'd5286: color_o = 12'b000011110000;
		13'd5287: color_o = 12'b000011110000;
		13'd5288: color_o = 12'b000011110000;
		13'd5289: color_o = 12'b000011110000;
		13'd5290: color_o = 12'b000011110000;
		13'd5291: color_o = 12'b000011110000;
		13'd5292: color_o = 12'b000011110000;
		13'd5293: color_o = 12'b000011110000;
		13'd5294: color_o = 12'b000011110000;
		13'd5295: color_o = 12'b000011110000;
		13'd5296: color_o = 12'b000011110000;
		13'd5297: color_o = 12'b000011110000;
		13'd5298: color_o = 12'b000011110000;
		13'd5299: color_o = 12'b000011110000;
		13'd5300: color_o = 12'b000011110000;
		13'd5301: color_o = 12'b000011110000;
		13'd5302: color_o = 12'b000011110000;
		13'd5303: color_o = 12'b000011110000;
		13'd5304: color_o = 12'b000011110000;
		13'd5305: color_o = 12'b000011110000;
		13'd5306: color_o = 12'b000011110000;
		13'd5307: color_o = 12'b000011110000;
		13'd5308: color_o = 12'b000011110000;
		13'd5309: color_o = 12'b000011110000;
		13'd5310: color_o = 12'b000011110000;
		13'd5311: color_o = 12'b000011110000;
		13'd5312: color_o = 12'b000011110000;
		13'd5313: color_o = 12'b000011110000;
		13'd5314: color_o = 12'b000011110000;
		13'd5315: color_o = 12'b000011110000;
		13'd5316: color_o = 12'b000011110000;
		13'd5317: color_o = 12'b000011110000;
		13'd5318: color_o = 12'b000000000000;
		13'd5319: color_o = 12'b000000000000;
		13'd5320: color_o = 12'b000000000000;
		13'd5321: color_o = 12'b000000000000;
		13'd5322: color_o = 12'b000000000000;
		13'd5323: color_o = 12'b000000000000;
		13'd5324: color_o = 12'b100000000000;
		13'd5325: color_o = 12'b100000000000;
		13'd5326: color_o = 12'b000000000000;
		13'd5327: color_o = 12'b000000000000;
		13'd5328: color_o = 12'b000000000000;
		13'd5329: color_o = 12'b100000000000;
		13'd5330: color_o = 12'b100000000000;
		13'd5331: color_o = 12'b000000000000;
		13'd5332: color_o = 12'b000000000000;
		13'd5333: color_o = 12'b000000000000;
		13'd5334: color_o = 12'b000000000000;
		13'd5335: color_o = 12'b000000000000;
		13'd5336: color_o = 12'b000000000000;
		13'd5337: color_o = 12'b000000000000;
		13'd5338: color_o = 12'b000000000000;
		13'd5339: color_o = 12'b000011110000;
		13'd5340: color_o = 12'b000011110000;
		13'd5341: color_o = 12'b000011110000;
		13'd5342: color_o = 12'b000011110000;
		13'd5343: color_o = 12'b000011110000;
		13'd5344: color_o = 12'b000011110000;
		13'd5345: color_o = 12'b000011110000;
		13'd5346: color_o = 12'b000011110000;
		13'd5347: color_o = 12'b000011110000;
		13'd5348: color_o = 12'b000011110000;
		13'd5349: color_o = 12'b000011110000;
		13'd5350: color_o = 12'b000011110000;
		13'd5351: color_o = 12'b000011110000;
		13'd5352: color_o = 12'b000011110000;
		13'd5353: color_o = 12'b000011110000;
		13'd5354: color_o = 12'b000011110000;
		13'd5355: color_o = 12'b000011110000;
		13'd5356: color_o = 12'b000011110000;
		13'd5357: color_o = 12'b000011110000;
		13'd5358: color_o = 12'b000011110000;
		13'd5359: color_o = 12'b000011110000;
		13'd5360: color_o = 12'b000011110000;
		13'd5361: color_o = 12'b000011110000;
		13'd5362: color_o = 12'b000011110000;
		13'd5363: color_o = 12'b000011110000;
		13'd5364: color_o = 12'b000011110000;
		13'd5365: color_o = 12'b000011110000;
		13'd5366: color_o = 12'b000011110000;
		13'd5367: color_o = 12'b000011110000;
		13'd5368: color_o = 12'b000011110000;
		13'd5369: color_o = 12'b000011110000;
		13'd5370: color_o = 12'b000011110000;
		13'd5371: color_o = 12'b000011110000;
		13'd5372: color_o = 12'b000011110000;
		13'd5373: color_o = 12'b000011110000;
		13'd5374: color_o = 12'b000011110000;
		13'd5375: color_o = 12'b000011110000;
		13'd5376: color_o = 12'b000011110000;
		13'd5377: color_o = 12'b000011110000;
		13'd5378: color_o = 12'b000011110000;
		13'd5379: color_o = 12'b000011110000;
		13'd5380: color_o = 12'b000011110000;
		13'd5381: color_o = 12'b000011110000;
		13'd5382: color_o = 12'b000011110000;
		13'd5383: color_o = 12'b000011110000;
		13'd5384: color_o = 12'b000011110000;
		13'd5385: color_o = 12'b000011110000;
		13'd5386: color_o = 12'b000011110000;
		13'd5387: color_o = 12'b000011110000;
		13'd5388: color_o = 12'b000011110000;
		13'd5389: color_o = 12'b000011110000;
		13'd5390: color_o = 12'b000011110000;
		13'd5391: color_o = 12'b000011110000;
		13'd5392: color_o = 12'b000011110000;
		13'd5393: color_o = 12'b000011110000;
		13'd5394: color_o = 12'b000011110000;
		13'd5395: color_o = 12'b000011110000;
		13'd5396: color_o = 12'b000011110000;
		13'd5397: color_o = 12'b000011110000;
		13'd5398: color_o = 12'b000011110000;
		13'd5399: color_o = 12'b000011110000;
		13'd5400: color_o = 12'b000011110000;
		13'd5401: color_o = 12'b000011110000;
		13'd5402: color_o = 12'b000011110000;
		13'd5403: color_o = 12'b000011110000;
		13'd5404: color_o = 12'b000011110000;
		13'd5405: color_o = 12'b000011110000;
		13'd5406: color_o = 12'b000011110000;
		13'd5407: color_o = 12'b000011110000;
		13'd5408: color_o = 12'b000011110000;
		13'd5409: color_o = 12'b000011110000;
		13'd5410: color_o = 12'b000011110000;
		13'd5411: color_o = 12'b000011110000;
		13'd5412: color_o = 12'b000011110000;
		13'd5413: color_o = 12'b000011110000;
		13'd5414: color_o = 12'b000011110000;
		13'd5415: color_o = 12'b000011110000;
		13'd5416: color_o = 12'b000011110000;
		13'd5417: color_o = 12'b000011110000;
		13'd5418: color_o = 12'b000011110000;
		13'd5419: color_o = 12'b000011110000;
		13'd5420: color_o = 12'b000011110000;
		13'd5421: color_o = 12'b000011110000;
		13'd5422: color_o = 12'b000011110000;
		13'd5423: color_o = 12'b000011110000;
		13'd5424: color_o = 12'b000011110000;
		13'd5425: color_o = 12'b000011110000;
		13'd5426: color_o = 12'b000011110000;
		13'd5427: color_o = 12'b000011110000;
		13'd5428: color_o = 12'b000011110000;
		13'd5429: color_o = 12'b000011110000;
		13'd5430: color_o = 12'b000011110000;
		13'd5431: color_o = 12'b000011110000;
		13'd5432: color_o = 12'b000011110000;
		13'd5433: color_o = 12'b000011110000;
		13'd5434: color_o = 12'b000011110000;
		13'd5435: color_o = 12'b000011110000;
		13'd5436: color_o = 12'b000011110000;
		13'd5437: color_o = 12'b000011110000;
		13'd5438: color_o = 12'b000011110000;
		13'd5439: color_o = 12'b000011110000;
		13'd5440: color_o = 12'b000011110000;
		13'd5441: color_o = 12'b000011110000;
		13'd5442: color_o = 12'b000011110000;
		13'd5443: color_o = 12'b000011110000;
		13'd5444: color_o = 12'b000011110000;
		13'd5445: color_o = 12'b000011110000;
		13'd5446: color_o = 12'b000011110000;
		13'd5447: color_o = 12'b000011110000;
		13'd5448: color_o = 12'b000011110000;
		13'd5449: color_o = 12'b000011110000;
		13'd5450: color_o = 12'b000011110000;
		13'd5451: color_o = 12'b000011110000;
		13'd5452: color_o = 12'b000011110000;
		13'd5453: color_o = 12'b000011110000;
		13'd5454: color_o = 12'b000011110000;
		13'd5455: color_o = 12'b000011110000;
		13'd5456: color_o = 12'b000011110000;
		13'd5457: color_o = 12'b000011110000;
		13'd5458: color_o = 12'b000011110000;
		13'd5459: color_o = 12'b000011110000;
		13'd5460: color_o = 12'b000011110000;
		13'd5461: color_o = 12'b000011110000;
		13'd5462: color_o = 12'b000011110000;
		13'd5463: color_o = 12'b000011110000;
		13'd5464: color_o = 12'b000011110000;
		13'd5465: color_o = 12'b000011110000;
		13'd5466: color_o = 12'b000011110000;
		13'd5467: color_o = 12'b000011110000;
		13'd5468: color_o = 12'b000011110000;
		13'd5469: color_o = 12'b000011110000;
		13'd5470: color_o = 12'b000011110000;
		13'd5471: color_o = 12'b000011110000;
		13'd5472: color_o = 12'b000011110000;
		13'd5473: color_o = 12'b000011110000;
		13'd5474: color_o = 12'b000011110000;
		13'd5475: color_o = 12'b000011110000;
		13'd5476: color_o = 12'b000011110000;
		13'd5477: color_o = 12'b000011110000;
		13'd5478: color_o = 12'b000011110000;
		13'd5479: color_o = 12'b000011110000;
		13'd5480: color_o = 12'b000011110000;
		13'd5481: color_o = 12'b000011110000;
		13'd5482: color_o = 12'b000011110000;
		13'd5483: color_o = 12'b000011110000;
		13'd5484: color_o = 12'b000011110000;
		13'd5485: color_o = 12'b000011110000;
		13'd5486: color_o = 12'b000011110000;
		13'd5487: color_o = 12'b000011110000;
		13'd5488: color_o = 12'b000011110000;
		13'd5489: color_o = 12'b000011110000;
		13'd5490: color_o = 12'b000011110000;
		13'd5491: color_o = 12'b000011110000;
		13'd5492: color_o = 12'b000011110000;
		13'd5493: color_o = 12'b000011110000;
		13'd5494: color_o = 12'b000011110000;
		13'd5495: color_o = 12'b000011110000;
		13'd5496: color_o = 12'b000011110000;
		13'd5497: color_o = 12'b000011110000;
		13'd5498: color_o = 12'b000011110000;
		13'd5499: color_o = 12'b000011110000;
		13'd5500: color_o = 12'b000011110000;
		13'd5501: color_o = 12'b000011110000;
		13'd5502: color_o = 12'b000011110000;
		13'd5503: color_o = 12'b000011110000;
		13'd5504: color_o = 12'b000011110000;
		13'd5505: color_o = 12'b000011110000;
		13'd5506: color_o = 12'b000011110000;
		13'd5507: color_o = 12'b000011110000;
		13'd5508: color_o = 12'b000011110000;
		13'd5509: color_o = 12'b000011110000;
		13'd5510: color_o = 12'b000011110000;
		13'd5511: color_o = 12'b000011110000;
		13'd5512: color_o = 12'b000011110000;
		13'd5513: color_o = 12'b000011110000;
		13'd5514: color_o = 12'b000011110000;
		13'd5515: color_o = 12'b000011110000;
		13'd5516: color_o = 12'b000011110000;
		13'd5517: color_o = 12'b000011110000;
		13'd5518: color_o = 12'b000011110000;
		13'd5519: color_o = 12'b000011110000;
		13'd5520: color_o = 12'b000011110000;
		13'd5521: color_o = 12'b000011110000;
		13'd5522: color_o = 12'b000011110000;
		13'd5523: color_o = 12'b000011110000;
		13'd5524: color_o = 12'b000011110000;
		13'd5525: color_o = 12'b000011110000;
		13'd5526: color_o = 12'b000011110000;
		13'd5527: color_o = 12'b000011110000;
		13'd5528: color_o = 12'b000011110000;
		13'd5529: color_o = 12'b000011110000;
		13'd5530: color_o = 12'b000011110000;
		13'd5531: color_o = 12'b000011110000;
		13'd5532: color_o = 12'b000011110000;
		13'd5533: color_o = 12'b000011110000;
		13'd5534: color_o = 12'b000011110000;
		13'd5535: color_o = 12'b000011110000;
		13'd5536: color_o = 12'b000011110000;
		13'd5537: color_o = 12'b000011110000;
		13'd5538: color_o = 12'b000011110000;
		13'd5539: color_o = 12'b000011110000;
		13'd5540: color_o = 12'b000011110000;
		13'd5541: color_o = 12'b000011110000;
		13'd5542: color_o = 12'b000011110000;
		13'd5543: color_o = 12'b000011110000;
		13'd5544: color_o = 12'b000011110000;
		13'd5545: color_o = 12'b000011110000;
		13'd5546: color_o = 12'b000011110000;
		13'd5547: color_o = 12'b000011110000;
		13'd5548: color_o = 12'b000011110000;
		13'd5549: color_o = 12'b000011110000;
		13'd5550: color_o = 12'b000011110000;
		13'd5551: color_o = 12'b000011110000;
		13'd5552: color_o = 12'b000011110000;
		13'd5553: color_o = 12'b000011110000;
		13'd5554: color_o = 12'b000011110000;
		13'd5555: color_o = 12'b000011110000;
		13'd5556: color_o = 12'b000011110000;
		13'd5557: color_o = 12'b000011110000;
		13'd5558: color_o = 12'b000011110000;
		13'd5559: color_o = 12'b000011110000;
		13'd5560: color_o = 12'b000011110000;
		13'd5561: color_o = 12'b000011110000;
		13'd5562: color_o = 12'b000011110000;
		13'd5563: color_o = 12'b000011110000;
		13'd5564: color_o = 12'b000011110000;
		13'd5565: color_o = 12'b000011110000;
		13'd5566: color_o = 12'b000011110000;
		13'd5567: color_o = 12'b000011110000;
		13'd5568: color_o = 12'b000011110000;
		13'd5569: color_o = 12'b000011110000;
		13'd5570: color_o = 12'b000011110000;
		13'd5571: color_o = 12'b000011110000;
		13'd5572: color_o = 12'b000011110000;
		13'd5573: color_o = 12'b000011110000;
		13'd5574: color_o = 12'b000011110000;
		13'd5575: color_o = 12'b000011110000;
		13'd5576: color_o = 12'b000011110000;
		13'd5577: color_o = 12'b000011110000;
		13'd5578: color_o = 12'b000011110000;
		13'd5579: color_o = 12'b000011110000;
		13'd5580: color_o = 12'b000011110000;
		13'd5581: color_o = 12'b000011110000;
		13'd5582: color_o = 12'b000011110000;
		13'd5583: color_o = 12'b000011110000;
		13'd5584: color_o = 12'b000011110000;
		13'd5585: color_o = 12'b000011110000;
		13'd5586: color_o = 12'b000011110000;
		13'd5587: color_o = 12'b000011110000;
		13'd5588: color_o = 12'b000011110000;
		13'd5589: color_o = 12'b000011110000;
		13'd5590: color_o = 12'b000011110000;
		13'd5591: color_o = 12'b000011110000;
		13'd5592: color_o = 12'b000011110000;
		13'd5593: color_o = 12'b000011110000;
		13'd5594: color_o = 12'b000011110000;
		13'd5595: color_o = 12'b000011110000;
		13'd5596: color_o = 12'b000011110000;
		13'd5597: color_o = 12'b000011110000;
		13'd5598: color_o = 12'b000011110000;
		13'd5599: color_o = 12'b000011110000;
		13'd5600: color_o = 12'b000011110000;
		13'd5601: color_o = 12'b000011110000;
		13'd5602: color_o = 12'b000011110000;
		13'd5603: color_o = 12'b000011110000;
		13'd5604: color_o = 12'b000011110000;
		13'd5605: color_o = 12'b000011110000;
		13'd5606: color_o = 12'b000011110000;
		13'd5607: color_o = 12'b000011110000;
		13'd5608: color_o = 12'b000011110000;
		13'd5609: color_o = 12'b000011110000;
		13'd5610: color_o = 12'b000011110000;
		13'd5611: color_o = 12'b000011110000;
		13'd5612: color_o = 12'b000011110000;
		13'd5613: color_o = 12'b000011110000;
		13'd5614: color_o = 12'b000011110000;
		13'd5615: color_o = 12'b000011110000;
		13'd5616: color_o = 12'b000011110000;
		13'd5617: color_o = 12'b000011110000;
		13'd5618: color_o = 12'b000011110000;
		13'd5619: color_o = 12'b000011110000;
		13'd5620: color_o = 12'b000011110000;
		13'd5621: color_o = 12'b000011110000;
		13'd5622: color_o = 12'b000011110000;
		13'd5623: color_o = 12'b000011110000;
		13'd5624: color_o = 12'b000011110000;
		13'd5625: color_o = 12'b000011110000;
		13'd5626: color_o = 12'b000011110000;
		13'd5627: color_o = 12'b000011110000;
		13'd5628: color_o = 12'b000011110000;
		13'd5629: color_o = 12'b000011110000;
		13'd5630: color_o = 12'b000011110000;
		13'd5631: color_o = 12'b000011110000;

        default: color_o = 12'h000;
    endcase       
    
endmodule
